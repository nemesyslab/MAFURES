//   Engineer aydin emre guzel
//   04/09/2016 19:15:12
`timescale 1 ns / 1 ps
module test_v1
	#( parameter BitWidth = 32 )
	(
	input rst,
	input [BitWidth-1:0] u_S1,
	input [BitWidth-1:0] u_S0,
	input [BitWidth-1:0] v_S1,
	input [BitWidth-1:0] v_S0,
	input [BitWidth-1:0] w_S1,
	input [BitWidth-1:0] w_S0,
	input [BitWidth-1:0] p0,
	input [BitWidth-1:0] p2,
	input [BitWidth-1:0] p4,
	input [BitWidth-1:0] jj,
	input [BitWidth-1:0] u_S2,
	input [BitWidth-1:0] v_S2,
	input [BitWidth-1:0] w_S2,
	input [BitWidth-1:0] p1,
	input [BitWidth-1:0] p3,
	input [BitWidth-1:0] p5,
	input [BitWidth-1:0] ii,
	input [BitWidth-1:0] p0Prev,
	input [BitWidth-1:0] p2Prev,
	input [BitWidth-1:0] p4Prev,
	input [BitWidth-1:0] p1S_1,
	input [BitWidth-1:0] p3S_1,
	input [BitWidth-1:0] p5S_1,
	input [BitWidth-1:0] uS,
	input [BitWidth-1:0] vS,
	input [BitWidth-1:0] wS,
	input [BitWidth-1:0] u0S,
	input [BitWidth-1:0] v0S,
	input [BitWidth-1:0] I_xS,
	input [BitWidth-1:0] I_yS,
	input [BitWidth-1:0] I_tS,
	input [BitWidth-1:0] I_grad_sqrS,
	input [BitWidth-1:0] beta,
	output reg [BitWidth-1:0] p0Out,
	output reg [BitWidth-1:0] p2Out,
	output reg [BitWidth-1:0] p4Out,
	output reg [BitWidth-1:0] p1Out,
	output reg [BitWidth-1:0] p3Out,
	output reg [BitWidth-1:0] p5Out,
	output reg [BitWidth-1:0] uOut,
	output reg [BitWidth-1:0] vOut,
	output reg [BitWidth-1:0] wOut,
	output reg [BitWidth-1:0] u_Out,
	output reg [BitWidth-1:0] v_Out,
	output reg [BitWidth-1:0] w_Out,
	input clk
	);
	reg [3:0] state, stateNext;
	always@(*) begin
		if(rst)begin
			stateNext = 0;
		end else begin
			stateNext = state + 1;
			if(state == 9 )begin
				stateNext = 0;
			end
		end
	end
	always@(posedge clk) begin
		state <= stateNext;
	end
	localparam sub = 1;
	localparam add = 0;
	localparam lt = 1;
	localparam gt = 2;
	localparam m = 588;
	localparam n = 384;
	localparam carpan1 = 32'h3f000000;
	localparam carpan2 = 32'h3f000000;
	localparam cons0 = 32'h3e4ccccd;
	localparam cons5 = 32'h3f000000;
	localparam TAU = 32'h3ecccccd;
	localparam BETA = 32'h3dcccccd;
	localparam ZERO = 0;
	localparam ONE = 32'h3F800000;
	localparam TWO = 32'h40000000;
	localparam MINUSONE = 32'hBF800000;
	reg [BitWidth-1:0] reg000,reg000Next; reg [BitWidth-1:0] reg001,reg001Next; reg [BitWidth-1:0] reg002,reg002Next; reg [BitWidth-1:0] reg003,reg003Next; reg [BitWidth-1:0] reg004,reg004Next; reg [BitWidth-1:0] reg005,reg005Next; reg [BitWidth-1:0] reg006,reg006Next; reg [BitWidth-1:0] reg007,reg007Next; reg [BitWidth-1:0] reg008,reg008Next; reg [BitWidth-1:0] reg009,reg009Next; reg [BitWidth-1:0] reg010,reg010Next; reg [BitWidth-1:0] reg011,reg011Next; reg [BitWidth-1:0] reg012,reg012Next; reg [BitWidth-1:0] reg013,reg013Next; reg [BitWidth-1:0] reg014,reg014Next; reg [BitWidth-1:0] reg015,reg015Next; reg [BitWidth-1:0] reg016,reg016Next; reg [BitWidth-1:0] reg017,reg017Next; reg [BitWidth-1:0] reg018,reg018Next; reg [BitWidth-1:0] reg019,reg019Next; 
	reg [BitWidth-1:0] reg020,reg020Next; reg [BitWidth-1:0] reg021,reg021Next; reg [BitWidth-1:0] reg022,reg022Next; reg [BitWidth-1:0] reg023,reg023Next; reg [BitWidth-1:0] reg024,reg024Next; reg [BitWidth-1:0] reg025,reg025Next; reg [BitWidth-1:0] reg026,reg026Next; reg [BitWidth-1:0] reg027,reg027Next; reg [BitWidth-1:0] reg028,reg028Next; reg [BitWidth-1:0] reg029,reg029Next; reg [BitWidth-1:0] reg030,reg030Next; reg [BitWidth-1:0] reg031,reg031Next; reg [BitWidth-1:0] reg032,reg032Next; reg [BitWidth-1:0] reg033,reg033Next; reg [BitWidth-1:0] reg034,reg034Next; reg [BitWidth-1:0] reg035,reg035Next; reg [BitWidth-1:0] reg036,reg036Next; reg [BitWidth-1:0] reg037,reg037Next; reg [BitWidth-1:0] reg038,reg038Next; reg [BitWidth-1:0] reg039,reg039Next; 
	reg [BitWidth-1:0] reg040,reg040Next; reg [BitWidth-1:0] reg041,reg041Next; reg [BitWidth-1:0] reg042,reg042Next; reg [BitWidth-1:0] reg043,reg043Next; reg [BitWidth-1:0] reg044,reg044Next; reg [BitWidth-1:0] reg045,reg045Next; reg [BitWidth-1:0] reg046,reg046Next; reg [BitWidth-1:0] reg047,reg047Next; reg [BitWidth-1:0] reg048,reg048Next; reg [BitWidth-1:0] reg049,reg049Next; reg [BitWidth-1:0] reg050,reg050Next; reg [BitWidth-1:0] reg051,reg051Next; reg [BitWidth-1:0] reg052,reg052Next; reg [BitWidth-1:0] reg053,reg053Next; reg [BitWidth-1:0] reg054,reg054Next; reg [BitWidth-1:0] reg055,reg055Next; reg [BitWidth-1:0] reg056,reg056Next; reg [BitWidth-1:0] reg057,reg057Next; reg [BitWidth-1:0] reg058,reg058Next; reg [BitWidth-1:0] reg059,reg059Next; 
	reg [BitWidth-1:0] reg060,reg060Next; reg [BitWidth-1:0] reg061,reg061Next; reg [BitWidth-1:0] reg062,reg062Next; reg [BitWidth-1:0] reg063,reg063Next; reg [BitWidth-1:0] reg064,reg064Next; reg [BitWidth-1:0] reg065,reg065Next; reg [BitWidth-1:0] reg066,reg066Next; reg [BitWidth-1:0] reg067,reg067Next; reg [BitWidth-1:0] reg068,reg068Next; reg [BitWidth-1:0] reg069,reg069Next; reg [BitWidth-1:0] reg070,reg070Next; reg [BitWidth-1:0] reg071,reg071Next; reg [BitWidth-1:0] reg072,reg072Next; reg [BitWidth-1:0] reg073,reg073Next; reg [BitWidth-1:0] reg074,reg074Next; reg [BitWidth-1:0] reg075,reg075Next; reg [BitWidth-1:0] reg076,reg076Next; reg [BitWidth-1:0] reg077,reg077Next; reg [BitWidth-1:0] reg078,reg078Next; reg [BitWidth-1:0] reg079,reg079Next; 
	reg [BitWidth-1:0] reg080,reg080Next; reg [BitWidth-1:0] reg081,reg081Next; reg [BitWidth-1:0] reg082,reg082Next; reg [BitWidth-1:0] reg083,reg083Next; reg [BitWidth-1:0] reg084,reg084Next; reg [BitWidth-1:0] reg085,reg085Next; reg [BitWidth-1:0] reg086,reg086Next; reg [BitWidth-1:0] reg087,reg087Next; reg [BitWidth-1:0] reg088,reg088Next; reg [BitWidth-1:0] reg089,reg089Next; reg [BitWidth-1:0] reg090,reg090Next; reg [BitWidth-1:0] reg091,reg091Next; reg [BitWidth-1:0] reg092,reg092Next; reg [BitWidth-1:0] reg093,reg093Next; reg [BitWidth-1:0] reg094,reg094Next; reg [BitWidth-1:0] reg095,reg095Next; reg [BitWidth-1:0] reg096,reg096Next; reg [BitWidth-1:0] reg097,reg097Next; reg [BitWidth-1:0] reg098,reg098Next; reg [BitWidth-1:0] reg099,reg099Next; 
	reg [BitWidth-1:0] reg100,reg100Next; reg [BitWidth-1:0] reg101,reg101Next; reg [BitWidth-1:0] reg102,reg102Next; reg [BitWidth-1:0] reg103,reg103Next; reg [BitWidth-1:0] reg104,reg104Next; reg [BitWidth-1:0] reg105,reg105Next; reg [BitWidth-1:0] reg106,reg106Next; reg [BitWidth-1:0] reg107,reg107Next; reg [BitWidth-1:0] reg108,reg108Next; reg [BitWidth-1:0] reg109,reg109Next; reg [BitWidth-1:0] reg110,reg110Next; reg [BitWidth-1:0] reg111,reg111Next; reg [BitWidth-1:0] reg112,reg112Next; reg [BitWidth-1:0] reg113,reg113Next; reg [BitWidth-1:0] reg114,reg114Next; reg [BitWidth-1:0] reg115,reg115Next; reg [BitWidth-1:0] reg116,reg116Next; reg [BitWidth-1:0] reg117,reg117Next; reg [BitWidth-1:0] reg118,reg118Next; reg [BitWidth-1:0] reg119,reg119Next; 
	reg [BitWidth-1:0] reg120,reg120Next; reg [BitWidth-1:0] reg121,reg121Next; reg [BitWidth-1:0] reg122,reg122Next; reg [BitWidth-1:0] reg123,reg123Next; reg [BitWidth-1:0] reg124,reg124Next; reg [BitWidth-1:0] reg125,reg125Next; reg [BitWidth-1:0] reg126,reg126Next; reg [BitWidth-1:0] reg127,reg127Next; reg [BitWidth-1:0] reg128,reg128Next; reg [BitWidth-1:0] reg129,reg129Next; reg [BitWidth-1:0] reg130,reg130Next; reg [BitWidth-1:0] reg131,reg131Next; reg [BitWidth-1:0] reg132,reg132Next; reg [BitWidth-1:0] reg133,reg133Next; reg [BitWidth-1:0] reg134,reg134Next; reg [BitWidth-1:0] reg135,reg135Next; reg [BitWidth-1:0] reg136,reg136Next; reg [BitWidth-1:0] reg137,reg137Next; reg [BitWidth-1:0] reg138,reg138Next; reg [BitWidth-1:0] reg139,reg139Next; 
	reg [BitWidth-1:0] reg140,reg140Next; reg [BitWidth-1:0] reg141,reg141Next; reg [BitWidth-1:0] reg142,reg142Next; reg [BitWidth-1:0] reg143,reg143Next; reg [BitWidth-1:0] reg144,reg144Next; reg [BitWidth-1:0] reg145,reg145Next; reg [BitWidth-1:0] reg146,reg146Next; reg [BitWidth-1:0] reg147,reg147Next; reg [BitWidth-1:0] reg148,reg148Next; reg [BitWidth-1:0] reg149,reg149Next; reg [BitWidth-1:0] reg150,reg150Next; reg [BitWidth-1:0] reg151,reg151Next; reg [BitWidth-1:0] reg152,reg152Next; reg [BitWidth-1:0] reg153,reg153Next; reg [BitWidth-1:0] reg154,reg154Next; reg [BitWidth-1:0] reg155,reg155Next; reg [BitWidth-1:0] reg156,reg156Next; reg [BitWidth-1:0] reg157,reg157Next; reg [BitWidth-1:0] reg158,reg158Next; reg [BitWidth-1:0] reg159,reg159Next; 
	reg [BitWidth-1:0] reg160,reg160Next; reg [BitWidth-1:0] reg161,reg161Next; reg [BitWidth-1:0] reg162,reg162Next; reg [BitWidth-1:0] reg163,reg163Next; reg [BitWidth-1:0] reg164,reg164Next; reg [BitWidth-1:0] reg165,reg165Next; reg [BitWidth-1:0] reg166,reg166Next; reg [BitWidth-1:0] reg167,reg167Next; reg [BitWidth-1:0] reg168,reg168Next; reg [BitWidth-1:0] reg169,reg169Next; reg [BitWidth-1:0] reg170,reg170Next; reg [BitWidth-1:0] reg171,reg171Next; reg [BitWidth-1:0] reg172,reg172Next; reg [BitWidth-1:0] reg173,reg173Next; reg [BitWidth-1:0] reg174,reg174Next; reg [BitWidth-1:0] reg175,reg175Next; reg [BitWidth-1:0] reg176,reg176Next; reg [BitWidth-1:0] reg177,reg177Next; reg [BitWidth-1:0] reg178,reg178Next; reg [BitWidth-1:0] reg179,reg179Next; 
	reg [BitWidth-1:0] reg180,reg180Next; reg [BitWidth-1:0] reg181,reg181Next; reg [BitWidth-1:0] reg182,reg182Next; reg [BitWidth-1:0] reg183,reg183Next; reg [BitWidth-1:0] reg184,reg184Next; reg [BitWidth-1:0] reg185,reg185Next; reg [BitWidth-1:0] reg186,reg186Next; reg [BitWidth-1:0] reg187,reg187Next; reg [BitWidth-1:0] reg188,reg188Next; reg [BitWidth-1:0] reg189,reg189Next; reg [BitWidth-1:0] reg190,reg190Next; reg [BitWidth-1:0] reg191,reg191Next; reg [BitWidth-1:0] reg192,reg192Next; reg [BitWidth-1:0] reg193,reg193Next; reg [BitWidth-1:0] reg194,reg194Next; reg [BitWidth-1:0] reg195,reg195Next; reg [BitWidth-1:0] reg196,reg196Next; reg [BitWidth-1:0] reg197,reg197Next; reg [BitWidth-1:0] reg198,reg198Next; reg [BitWidth-1:0] reg199,reg199Next; 
	reg [BitWidth-1:0] reg200,reg200Next; reg [BitWidth-1:0] reg201,reg201Next; reg [BitWidth-1:0] reg202,reg202Next; reg [BitWidth-1:0] reg203,reg203Next; reg [BitWidth-1:0] reg204,reg204Next; reg [BitWidth-1:0] reg205,reg205Next; reg [BitWidth-1:0] reg206,reg206Next; reg [BitWidth-1:0] reg207,reg207Next; reg [BitWidth-1:0] reg208,reg208Next; reg [BitWidth-1:0] reg209,reg209Next; reg [BitWidth-1:0] reg210,reg210Next; reg [BitWidth-1:0] reg211,reg211Next; reg [BitWidth-1:0] reg212,reg212Next; reg [BitWidth-1:0] reg213,reg213Next; reg [BitWidth-1:0] reg214,reg214Next; reg [BitWidth-1:0] reg215,reg215Next; reg [BitWidth-1:0] reg216,reg216Next; reg [BitWidth-1:0] reg217,reg217Next; reg [BitWidth-1:0] reg218,reg218Next; reg [BitWidth-1:0] reg219,reg219Next; 
	reg [BitWidth-1:0] reg220,reg220Next; reg [BitWidth-1:0] reg221,reg221Next; reg [BitWidth-1:0] reg222,reg222Next; reg [BitWidth-1:0] reg223,reg223Next; reg [BitWidth-1:0] reg224,reg224Next; reg [BitWidth-1:0] reg225,reg225Next; reg [BitWidth-1:0] reg226,reg226Next; reg [BitWidth-1:0] reg227,reg227Next; reg [BitWidth-1:0] reg228,reg228Next; reg [BitWidth-1:0] reg229,reg229Next; reg [BitWidth-1:0] reg230,reg230Next; reg [BitWidth-1:0] reg231,reg231Next; reg [BitWidth-1:0] reg232,reg232Next; reg [BitWidth-1:0] reg233,reg233Next; reg [BitWidth-1:0] reg234,reg234Next; reg [BitWidth-1:0] reg235,reg235Next; reg [BitWidth-1:0] reg236,reg236Next; reg [BitWidth-1:0] reg237,reg237Next; reg [BitWidth-1:0] reg238,reg238Next; reg [BitWidth-1:0] reg239,reg239Next; 
	reg [BitWidth-1:0] reg240,reg240Next; reg [BitWidth-1:0] reg241,reg241Next; reg [BitWidth-1:0] reg242,reg242Next; reg [BitWidth-1:0] reg243,reg243Next; reg [BitWidth-1:0] reg244,reg244Next; reg [BitWidth-1:0] reg245,reg245Next; reg [BitWidth-1:0] reg246,reg246Next; reg [BitWidth-1:0] reg247,reg247Next; reg [BitWidth-1:0] reg248,reg248Next; reg [BitWidth-1:0] reg249,reg249Next; reg [BitWidth-1:0] reg250,reg250Next; reg [BitWidth-1:0] reg251,reg251Next; reg [BitWidth-1:0] reg252,reg252Next; reg [BitWidth-1:0] reg253,reg253Next; reg [BitWidth-1:0] reg254,reg254Next; reg [BitWidth-1:0] reg255,reg255Next; reg [BitWidth-1:0] reg256,reg256Next; reg [BitWidth-1:0] reg257,reg257Next; reg [BitWidth-1:0] reg258,reg258Next; reg [BitWidth-1:0] reg259,reg259Next; 
	reg [BitWidth-1:0] reg260,reg260Next; reg [BitWidth-1:0] reg261,reg261Next; reg [BitWidth-1:0] reg262,reg262Next; reg [BitWidth-1:0] reg263,reg263Next; reg [BitWidth-1:0] reg264,reg264Next; reg [BitWidth-1:0] reg265,reg265Next; reg [BitWidth-1:0] reg266,reg266Next; reg [BitWidth-1:0] reg267,reg267Next; reg [BitWidth-1:0] reg268,reg268Next; reg [BitWidth-1:0] reg269,reg269Next; reg [BitWidth-1:0] reg270,reg270Next; reg [BitWidth-1:0] reg271,reg271Next; reg [BitWidth-1:0] reg272,reg272Next; reg [BitWidth-1:0] reg273,reg273Next; reg [BitWidth-1:0] reg274,reg274Next; reg [BitWidth-1:0] reg275,reg275Next; reg [BitWidth-1:0] reg276,reg276Next; reg [BitWidth-1:0] reg277,reg277Next; reg [BitWidth-1:0] reg278,reg278Next; reg [BitWidth-1:0] reg279,reg279Next; 
	reg [BitWidth-1:0] reg280,reg280Next; reg [BitWidth-1:0] reg281,reg281Next; reg [BitWidth-1:0] reg282,reg282Next; reg [BitWidth-1:0] reg283,reg283Next; reg [BitWidth-1:0] reg284,reg284Next; reg [BitWidth-1:0] reg285,reg285Next; reg [BitWidth-1:0] reg286,reg286Next; reg [BitWidth-1:0] reg287,reg287Next; reg [BitWidth-1:0] reg288,reg288Next; reg [BitWidth-1:0] reg289,reg289Next; reg [BitWidth-1:0] reg290,reg290Next; reg [BitWidth-1:0] reg291,reg291Next; reg [BitWidth-1:0] reg292,reg292Next; reg [BitWidth-1:0] reg293,reg293Next; reg [BitWidth-1:0] reg294,reg294Next; reg [BitWidth-1:0] reg295,reg295Next; reg [BitWidth-1:0] reg296,reg296Next; reg [BitWidth-1:0] reg297,reg297Next; reg [BitWidth-1:0] reg298,reg298Next; reg [BitWidth-1:0] reg299,reg299Next; 
	reg [BitWidth-1:0] reg300,reg300Next; reg [BitWidth-1:0] reg301,reg301Next; reg [BitWidth-1:0] reg302,reg302Next; reg [BitWidth-1:0] reg303,reg303Next; reg [BitWidth-1:0] reg304,reg304Next; reg [BitWidth-1:0] reg305,reg305Next; reg [BitWidth-1:0] reg306,reg306Next; reg [BitWidth-1:0] reg307,reg307Next; reg [BitWidth-1:0] reg308,reg308Next; reg [BitWidth-1:0] reg309,reg309Next; reg [BitWidth-1:0] reg310,reg310Next; reg [BitWidth-1:0] reg311,reg311Next; reg [BitWidth-1:0] reg312,reg312Next; reg [BitWidth-1:0] reg313,reg313Next; reg [BitWidth-1:0] reg314,reg314Next; reg [BitWidth-1:0] reg315,reg315Next; reg [BitWidth-1:0] reg316,reg316Next; reg [BitWidth-1:0] reg317,reg317Next; reg [BitWidth-1:0] reg318,reg318Next; reg [BitWidth-1:0] reg319,reg319Next; 
	reg [BitWidth-1:0] reg320,reg320Next; reg [BitWidth-1:0] reg321,reg321Next; reg [BitWidth-1:0] reg322,reg322Next; reg [BitWidth-1:0] reg323,reg323Next; reg [BitWidth-1:0] reg324,reg324Next; reg [BitWidth-1:0] reg325,reg325Next; reg [BitWidth-1:0] reg326,reg326Next; reg [BitWidth-1:0] reg327,reg327Next; reg [BitWidth-1:0] reg328,reg328Next; reg [BitWidth-1:0] reg329,reg329Next; reg [BitWidth-1:0] reg330,reg330Next; reg [BitWidth-1:0] reg331,reg331Next; reg [BitWidth-1:0] reg332,reg332Next; reg [BitWidth-1:0] reg333,reg333Next; reg [BitWidth-1:0] reg334,reg334Next; reg [BitWidth-1:0] reg335,reg335Next; reg [BitWidth-1:0] reg336,reg336Next; reg [BitWidth-1:0] reg337,reg337Next; reg [BitWidth-1:0] reg338,reg338Next; reg [BitWidth-1:0] reg339,reg339Next; 
	reg [BitWidth-1:0] reg340,reg340Next; reg [BitWidth-1:0] reg341,reg341Next; reg [BitWidth-1:0] reg342,reg342Next; reg [BitWidth-1:0] reg343,reg343Next; reg [BitWidth-1:0] reg344,reg344Next; reg [BitWidth-1:0] reg345,reg345Next; reg [BitWidth-1:0] reg346,reg346Next; reg [BitWidth-1:0] reg347,reg347Next; reg [BitWidth-1:0] reg348,reg348Next; reg [BitWidth-1:0] reg349,reg349Next; reg [BitWidth-1:0] reg350,reg350Next; reg [BitWidth-1:0] reg351,reg351Next; reg [BitWidth-1:0] reg352,reg352Next; reg [BitWidth-1:0] reg353,reg353Next; reg [BitWidth-1:0] reg354,reg354Next; reg [BitWidth-1:0] reg355,reg355Next; reg [BitWidth-1:0] reg356,reg356Next; reg [BitWidth-1:0] reg357,reg357Next; reg [BitWidth-1:0] reg358,reg358Next; reg [BitWidth-1:0] reg359,reg359Next; 
	reg [BitWidth-1:0] reg360,reg360Next; reg [BitWidth-1:0] reg361,reg361Next; reg [BitWidth-1:0] reg362,reg362Next; reg [BitWidth-1:0] reg363,reg363Next; reg [BitWidth-1:0] reg364,reg364Next; reg [BitWidth-1:0] reg365,reg365Next; reg [BitWidth-1:0] reg366,reg366Next; reg [BitWidth-1:0] reg367,reg367Next; reg [BitWidth-1:0] reg368,reg368Next; reg [BitWidth-1:0] reg369,reg369Next; reg [BitWidth-1:0] reg370,reg370Next; reg [BitWidth-1:0] reg371,reg371Next; reg [BitWidth-1:0] reg372,reg372Next; reg [BitWidth-1:0] reg373,reg373Next; reg [BitWidth-1:0] reg374,reg374Next; reg [BitWidth-1:0] reg375,reg375Next; reg [BitWidth-1:0] reg376,reg376Next; reg [BitWidth-1:0] reg377,reg377Next; reg [BitWidth-1:0] reg378,reg378Next; reg [BitWidth-1:0] reg379,reg379Next; 
	reg [BitWidth-1:0] reg380,reg380Next; reg [BitWidth-1:0] reg381,reg381Next; reg [BitWidth-1:0] reg382,reg382Next; reg [BitWidth-1:0] reg383,reg383Next; reg [BitWidth-1:0] reg384,reg384Next; reg [BitWidth-1:0] reg385,reg385Next; reg [BitWidth-1:0] reg386,reg386Next; reg [BitWidth-1:0] reg387,reg387Next; reg [BitWidth-1:0] reg388,reg388Next; reg [BitWidth-1:0] reg389,reg389Next; reg [BitWidth-1:0] reg390,reg390Next; reg [BitWidth-1:0] reg391,reg391Next; reg [BitWidth-1:0] reg392,reg392Next; reg [BitWidth-1:0] reg393,reg393Next; reg [BitWidth-1:0] reg394,reg394Next; reg [BitWidth-1:0] reg395,reg395Next; reg [BitWidth-1:0] reg396,reg396Next; reg [BitWidth-1:0] reg397,reg397Next; reg [BitWidth-1:0] reg398,reg398Next; reg [BitWidth-1:0] reg399,reg399Next; 
	reg [BitWidth-1:0] reg400,reg400Next; reg [BitWidth-1:0] reg401,reg401Next; reg [BitWidth-1:0] reg402,reg402Next; reg [BitWidth-1:0] reg403,reg403Next; reg [BitWidth-1:0] reg404,reg404Next; reg [BitWidth-1:0] reg405,reg405Next; reg [BitWidth-1:0] reg406,reg406Next; reg [BitWidth-1:0] reg407,reg407Next; reg [BitWidth-1:0] reg408,reg408Next; reg [BitWidth-1:0] reg409,reg409Next; reg [BitWidth-1:0] reg410,reg410Next; reg [BitWidth-1:0] reg411,reg411Next; reg [BitWidth-1:0] reg412,reg412Next; reg [BitWidth-1:0] reg413,reg413Next; reg [BitWidth-1:0] reg414,reg414Next; reg [BitWidth-1:0] reg415,reg415Next; reg [BitWidth-1:0] reg416,reg416Next; reg [BitWidth-1:0] reg417,reg417Next; reg [BitWidth-1:0] reg418,reg418Next; reg [BitWidth-1:0] reg419,reg419Next; 
	reg [BitWidth-1:0] reg420,reg420Next; reg [BitWidth-1:0] reg421,reg421Next; reg [BitWidth-1:0] reg422,reg422Next; reg [BitWidth-1:0] reg423,reg423Next; reg [BitWidth-1:0] reg424,reg424Next; reg [BitWidth-1:0] reg425,reg425Next; reg [BitWidth-1:0] reg426,reg426Next; reg [BitWidth-1:0] reg427,reg427Next; reg [BitWidth-1:0] reg428,reg428Next; reg [BitWidth-1:0] reg429,reg429Next; reg [BitWidth-1:0] reg430,reg430Next; reg [BitWidth-1:0] reg431,reg431Next; reg [BitWidth-1:0] reg432,reg432Next; reg [BitWidth-1:0] reg433,reg433Next; reg [BitWidth-1:0] reg434,reg434Next; reg [BitWidth-1:0] reg435,reg435Next; reg [BitWidth-1:0] reg436,reg436Next; reg [BitWidth-1:0] reg437,reg437Next; reg [BitWidth-1:0] reg438,reg438Next; reg [BitWidth-1:0] reg439,reg439Next; 
	reg [BitWidth-1:0] reg440,reg440Next; reg [BitWidth-1:0] reg441,reg441Next; reg [BitWidth-1:0] reg442,reg442Next; reg [BitWidth-1:0] reg443,reg443Next; reg [BitWidth-1:0] reg444,reg444Next; reg [BitWidth-1:0] reg445,reg445Next; reg [BitWidth-1:0] reg446,reg446Next; reg [BitWidth-1:0] reg447,reg447Next; reg [BitWidth-1:0] reg448,reg448Next; reg [BitWidth-1:0] reg449,reg449Next; reg [BitWidth-1:0] reg450,reg450Next; reg [BitWidth-1:0] reg451,reg451Next; reg [BitWidth-1:0] reg452,reg452Next; reg [BitWidth-1:0] reg453,reg453Next; reg [BitWidth-1:0] reg454,reg454Next; reg [BitWidth-1:0] reg455,reg455Next; reg [BitWidth-1:0] reg456,reg456Next; reg [BitWidth-1:0] reg457,reg457Next; reg [BitWidth-1:0] reg458,reg458Next; reg [BitWidth-1:0] reg459,reg459Next; 
	reg [BitWidth-1:0] reg460,reg460Next; reg [BitWidth-1:0] reg461,reg461Next; reg [BitWidth-1:0] reg462,reg462Next; reg [BitWidth-1:0] reg463,reg463Next; reg [BitWidth-1:0] reg464,reg464Next; reg [BitWidth-1:0] reg465,reg465Next; reg [BitWidth-1:0] reg466,reg466Next; reg [BitWidth-1:0] reg467,reg467Next; reg [BitWidth-1:0] reg468,reg468Next; reg [BitWidth-1:0] reg469,reg469Next; reg [BitWidth-1:0] reg470,reg470Next; reg [BitWidth-1:0] reg471,reg471Next; reg [BitWidth-1:0] reg472,reg472Next; reg [BitWidth-1:0] reg473,reg473Next; reg [BitWidth-1:0] reg474,reg474Next; reg [BitWidth-1:0] reg475,reg475Next; reg [BitWidth-1:0] reg476,reg476Next; reg [BitWidth-1:0] reg477,reg477Next; reg [BitWidth-1:0] reg478,reg478Next; reg [BitWidth-1:0] reg479,reg479Next; 
	reg [BitWidth-1:0] reg480,reg480Next; reg [BitWidth-1:0] reg481,reg481Next; reg [BitWidth-1:0] reg482,reg482Next; reg [BitWidth-1:0] reg483,reg483Next; reg [BitWidth-1:0] reg484,reg484Next; reg [BitWidth-1:0] reg485,reg485Next; reg [BitWidth-1:0] reg486,reg486Next; reg [BitWidth-1:0] reg487,reg487Next; reg [BitWidth-1:0] reg488,reg488Next; reg [BitWidth-1:0] reg489,reg489Next; reg [BitWidth-1:0] reg490,reg490Next; reg [BitWidth-1:0] reg491,reg491Next; reg [BitWidth-1:0] reg492,reg492Next; reg [BitWidth-1:0] reg493,reg493Next; reg [BitWidth-1:0] reg494,reg494Next; reg [BitWidth-1:0] reg495,reg495Next; reg [BitWidth-1:0] reg496,reg496Next; reg [BitWidth-1:0] reg497,reg497Next; reg [BitWidth-1:0] reg498,reg498Next; reg [BitWidth-1:0] reg499,reg499Next; 
	reg [BitWidth-1:0] reg500,reg500Next; reg [BitWidth-1:0] reg501,reg501Next; reg [BitWidth-1:0] reg502,reg502Next; reg [BitWidth-1:0] reg503,reg503Next; reg [BitWidth-1:0] reg504,reg504Next; reg [BitWidth-1:0] reg505,reg505Next; reg [BitWidth-1:0] reg506,reg506Next; reg [BitWidth-1:0] reg507,reg507Next; reg [BitWidth-1:0] reg508,reg508Next; reg [BitWidth-1:0] reg509,reg509Next; reg [BitWidth-1:0] reg510,reg510Next; reg [BitWidth-1:0] reg511,reg511Next; reg [BitWidth-1:0] reg512,reg512Next; reg [BitWidth-1:0] reg513,reg513Next; reg [BitWidth-1:0] reg514,reg514Next; reg [BitWidth-1:0] reg515,reg515Next; reg [BitWidth-1:0] reg516,reg516Next; reg [BitWidth-1:0] reg517,reg517Next; reg [BitWidth-1:0] reg518,reg518Next; reg [BitWidth-1:0] reg519,reg519Next; 
	reg [BitWidth-1:0] reg520,reg520Next; reg [BitWidth-1:0] reg521,reg521Next; reg [BitWidth-1:0] reg522,reg522Next; reg [BitWidth-1:0] reg523,reg523Next; reg [BitWidth-1:0] reg524,reg524Next; reg [BitWidth-1:0] reg525,reg525Next; reg [BitWidth-1:0] reg526,reg526Next; reg [BitWidth-1:0] reg527,reg527Next; reg [BitWidth-1:0] reg528,reg528Next; reg [BitWidth-1:0] reg529,reg529Next; reg [BitWidth-1:0] reg530,reg530Next; reg [BitWidth-1:0] reg531,reg531Next; reg [BitWidth-1:0] reg532,reg532Next; reg [BitWidth-1:0] reg533,reg533Next; reg [BitWidth-1:0] reg534,reg534Next; reg [BitWidth-1:0] reg535,reg535Next; reg [BitWidth-1:0] reg536,reg536Next; reg [BitWidth-1:0] reg537,reg537Next; reg [BitWidth-1:0] reg538,reg538Next; reg [BitWidth-1:0] reg539,reg539Next; 
	reg [BitWidth-1:0] reg540,reg540Next; reg [BitWidth-1:0] reg541,reg541Next; reg [BitWidth-1:0] reg542,reg542Next; reg [BitWidth-1:0] reg543,reg543Next; reg [BitWidth-1:0] reg544,reg544Next; reg [BitWidth-1:0] reg545,reg545Next; reg [BitWidth-1:0] reg546,reg546Next; reg [BitWidth-1:0] reg547,reg547Next; reg [BitWidth-1:0] reg548,reg548Next; reg [BitWidth-1:0] reg549,reg549Next; reg [BitWidth-1:0] reg550,reg550Next; reg [BitWidth-1:0] reg551,reg551Next; reg [BitWidth-1:0] reg552,reg552Next; reg [BitWidth-1:0] reg553,reg553Next; reg [BitWidth-1:0] reg554,reg554Next; reg [BitWidth-1:0] reg555,reg555Next; reg [BitWidth-1:0] reg556,reg556Next; reg [BitWidth-1:0] reg557,reg557Next; reg [BitWidth-1:0] reg558,reg558Next; reg [BitWidth-1:0] reg559,reg559Next; 
	reg [BitWidth-1:0] reg560,reg560Next; reg [BitWidth-1:0] reg561,reg561Next; reg [BitWidth-1:0] reg562,reg562Next; reg [BitWidth-1:0] reg563,reg563Next; reg [BitWidth-1:0] reg564,reg564Next; reg [BitWidth-1:0] reg565,reg565Next; reg [BitWidth-1:0] reg566,reg566Next; reg [BitWidth-1:0] reg567,reg567Next; reg [BitWidth-1:0] reg568,reg568Next; reg [BitWidth-1:0] reg569,reg569Next; reg [BitWidth-1:0] reg570,reg570Next; reg [BitWidth-1:0] reg571,reg571Next; reg [BitWidth-1:0] reg572,reg572Next; reg [BitWidth-1:0] reg573,reg573Next; reg [BitWidth-1:0] reg574,reg574Next; reg [BitWidth-1:0] reg575,reg575Next; reg [BitWidth-1:0] reg576,reg576Next; reg [BitWidth-1:0] reg577,reg577Next; reg [BitWidth-1:0] reg578,reg578Next; reg [BitWidth-1:0] reg579,reg579Next; 
	reg [BitWidth-1:0] reg580,reg580Next; reg [BitWidth-1:0] reg581,reg581Next; reg [BitWidth-1:0] reg582,reg582Next; reg [BitWidth-1:0] reg583,reg583Next; reg [BitWidth-1:0] reg584,reg584Next; reg [BitWidth-1:0] reg585,reg585Next; reg [BitWidth-1:0] reg586,reg586Next; reg [BitWidth-1:0] reg587,reg587Next; reg [BitWidth-1:0] reg588,reg588Next; reg [BitWidth-1:0] reg589,reg589Next; reg [BitWidth-1:0] reg590,reg590Next; reg [BitWidth-1:0] reg591,reg591Next; reg [BitWidth-1:0] reg592,reg592Next; reg [BitWidth-1:0] reg593,reg593Next; reg [BitWidth-1:0] reg594,reg594Next; reg [BitWidth-1:0] reg595,reg595Next; reg [BitWidth-1:0] reg596,reg596Next; reg [BitWidth-1:0] reg597,reg597Next; reg [BitWidth-1:0] reg598,reg598Next; reg [BitWidth-1:0] reg599,reg599Next; 
	reg [BitWidth-1:0] reg600,reg600Next; reg [BitWidth-1:0] reg601,reg601Next; reg [BitWidth-1:0] reg602,reg602Next; reg [BitWidth-1:0] reg603,reg603Next; reg [BitWidth-1:0] reg604,reg604Next; reg [BitWidth-1:0] reg605,reg605Next; reg [BitWidth-1:0] reg606,reg606Next; reg [BitWidth-1:0] reg607,reg607Next; reg [BitWidth-1:0] reg608,reg608Next; reg [BitWidth-1:0] reg609,reg609Next; reg [BitWidth-1:0] reg610,reg610Next; reg [BitWidth-1:0] reg611,reg611Next; reg [BitWidth-1:0] reg612,reg612Next; reg [BitWidth-1:0] reg613,reg613Next; reg [BitWidth-1:0] reg614,reg614Next; reg [BitWidth-1:0] reg615,reg615Next; reg [BitWidth-1:0] reg616,reg616Next; reg [BitWidth-1:0] reg617,reg617Next; reg [BitWidth-1:0] reg618,reg618Next; reg [BitWidth-1:0] reg619,reg619Next; 
	reg [BitWidth-1:0] reg620,reg620Next; reg [BitWidth-1:0] reg621,reg621Next; reg [BitWidth-1:0] reg622,reg622Next; reg [BitWidth-1:0] reg623,reg623Next; reg [BitWidth-1:0] reg624,reg624Next; reg [BitWidth-1:0] reg625,reg625Next; reg [BitWidth-1:0] reg626,reg626Next; reg [BitWidth-1:0] reg627,reg627Next; reg [BitWidth-1:0] reg628,reg628Next; reg [BitWidth-1:0] reg629,reg629Next; reg [BitWidth-1:0] reg630,reg630Next; reg [BitWidth-1:0] reg631,reg631Next; reg [BitWidth-1:0] reg632,reg632Next; reg [BitWidth-1:0] reg633,reg633Next; reg [BitWidth-1:0] reg634,reg634Next; reg [BitWidth-1:0] reg635,reg635Next; reg [BitWidth-1:0] reg636,reg636Next; reg [BitWidth-1:0] reg637,reg637Next; reg [BitWidth-1:0] reg638,reg638Next; reg [BitWidth-1:0] reg639,reg639Next; 
	reg [BitWidth-1:0] reg640,reg640Next; reg [BitWidth-1:0] reg641,reg641Next; reg [BitWidth-1:0] reg642,reg642Next; reg [BitWidth-1:0] reg643,reg643Next; reg [BitWidth-1:0] reg644,reg644Next; reg [BitWidth-1:0] reg645,reg645Next; reg [BitWidth-1:0] reg646,reg646Next; reg [BitWidth-1:0] reg647,reg647Next; reg [BitWidth-1:0] reg648,reg648Next; reg [BitWidth-1:0] reg649,reg649Next; reg [BitWidth-1:0] reg650,reg650Next; reg [BitWidth-1:0] reg651,reg651Next; reg [BitWidth-1:0] reg652,reg652Next; reg [BitWidth-1:0] reg653,reg653Next; reg [BitWidth-1:0] reg654,reg654Next; reg [BitWidth-1:0] reg655,reg655Next; reg [BitWidth-1:0] reg656,reg656Next; reg [BitWidth-1:0] reg657,reg657Next; reg [BitWidth-1:0] reg658,reg658Next; reg [BitWidth-1:0] reg659,reg659Next; 
	reg [BitWidth-1:0] reg660,reg660Next; reg [BitWidth-1:0] reg661,reg661Next; reg [BitWidth-1:0] reg662,reg662Next; reg [BitWidth-1:0] reg663,reg663Next; reg [BitWidth-1:0] reg664,reg664Next; reg [BitWidth-1:0] reg665,reg665Next; reg [BitWidth-1:0] reg666,reg666Next; reg [BitWidth-1:0] reg667,reg667Next; reg [BitWidth-1:0] reg668,reg668Next; reg [BitWidth-1:0] reg669,reg669Next; reg [BitWidth-1:0] reg670,reg670Next; reg [BitWidth-1:0] reg671,reg671Next; reg [BitWidth-1:0] reg672,reg672Next; reg [BitWidth-1:0] reg673,reg673Next; reg [BitWidth-1:0] reg674,reg674Next; reg [BitWidth-1:0] reg675,reg675Next; reg [BitWidth-1:0] reg676,reg676Next; reg [BitWidth-1:0] reg677,reg677Next; reg [BitWidth-1:0] reg678,reg678Next; reg [BitWidth-1:0] reg679,reg679Next; 
	reg [BitWidth-1:0] reg680,reg680Next; reg [BitWidth-1:0] reg681,reg681Next; reg [BitWidth-1:0] reg682,reg682Next; reg [BitWidth-1:0] reg683,reg683Next; reg [BitWidth-1:0] reg684,reg684Next; reg [BitWidth-1:0] reg685,reg685Next; reg [BitWidth-1:0] reg686,reg686Next; reg [BitWidth-1:0] reg687,reg687Next; reg [BitWidth-1:0] reg688,reg688Next; reg [BitWidth-1:0] reg689,reg689Next; reg [BitWidth-1:0] reg690,reg690Next; reg [BitWidth-1:0] reg691,reg691Next; reg [BitWidth-1:0] reg692,reg692Next; reg [BitWidth-1:0] reg693,reg693Next; reg [BitWidth-1:0] reg694,reg694Next; reg [BitWidth-1:0] reg695,reg695Next; reg [BitWidth-1:0] reg696,reg696Next; reg [BitWidth-1:0] reg697,reg697Next; reg [BitWidth-1:0] reg698,reg698Next; reg [BitWidth-1:0] reg699,reg699Next; 
	reg [BitWidth-1:0] reg700,reg700Next; reg [BitWidth-1:0] reg701,reg701Next; reg [BitWidth-1:0] reg702,reg702Next; reg [BitWidth-1:0] reg703,reg703Next; reg [BitWidth-1:0] reg704,reg704Next; reg [BitWidth-1:0] reg705,reg705Next; reg [BitWidth-1:0] reg706,reg706Next; reg [BitWidth-1:0] reg707,reg707Next; reg [BitWidth-1:0] reg708,reg708Next; reg [BitWidth-1:0] reg709,reg709Next; reg [BitWidth-1:0] reg710,reg710Next; reg [BitWidth-1:0] reg711,reg711Next; reg [BitWidth-1:0] reg712,reg712Next; reg [BitWidth-1:0] reg713,reg713Next; reg [BitWidth-1:0] reg714,reg714Next; reg [BitWidth-1:0] reg715,reg715Next; reg [BitWidth-1:0] reg716,reg716Next; reg [BitWidth-1:0] reg717,reg717Next; reg [BitWidth-1:0] reg718,reg718Next; 
	reg [BitWidth-1:0] addsubIn0a, addsubIn0b;
	reg [BitWidth-1:0] addsubMod0Next; reg [BitWidth-1:0] addsubMod0;
	reg [BitWidth-1:0] addsubIn0aNext, addsubIn0bNext;
	wire [BitWidth-1:0] addsubOut0Next; reg [BitWidth-1:0] addsubOut0;
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp #(
		.ID(1),
		.NUM_STAGE(14),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp_U0(
		.clk(clk),
		.reset(rst),
		.din0(addsubIn0a),
		.din1(addsubIn0b),
		.opcode(addsubMod0),
		.ce(1'b1),
		.dout(addsubOut0Next)
	);
	reg [BitWidth-1:0] addsubIn1a, addsubIn1b;
	reg [BitWidth-1:0] addsubMod1Next; reg [BitWidth-1:0] addsubMod1;
	reg [BitWidth-1:0] addsubIn1aNext, addsubIn1bNext;
	wire [BitWidth-1:0] addsubOut1Next; reg [BitWidth-1:0] addsubOut1;
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp #(
		.ID(1),
		.NUM_STAGE(14),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp_U1(
		.clk(clk),
		.reset(rst),
		.din0(addsubIn1a),
		.din1(addsubIn1b),
		.opcode(addsubMod1),
		.ce(1'b1),
		.dout(addsubOut1Next)
	);
	reg [BitWidth-1:0] addsubIn2a, addsubIn2b;
	reg [BitWidth-1:0] addsubMod2Next; reg [BitWidth-1:0] addsubMod2;
	reg [BitWidth-1:0] addsubIn2aNext, addsubIn2bNext;
	wire [BitWidth-1:0] addsubOut2Next; reg [BitWidth-1:0] addsubOut2;
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp #(
		.ID(1),
		.NUM_STAGE(14),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp_U2(
		.clk(clk),
		.reset(rst),
		.din0(addsubIn2a),
		.din1(addsubIn2b),
		.opcode(addsubMod2),
		.ce(1'b1),
		.dout(addsubOut2Next)
	);
	reg [BitWidth-1:0] addsubIn3a, addsubIn3b;
	reg [BitWidth-1:0] addsubMod3Next; reg [BitWidth-1:0] addsubMod3;
	reg [BitWidth-1:0] addsubIn3aNext, addsubIn3bNext;
	wire [BitWidth-1:0] addsubOut3Next; reg [BitWidth-1:0] addsubOut3;
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp #(
		.ID(1),
		.NUM_STAGE(14),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_faddfsub_32ns_32ns_32_14_no_dsp_U3(
		.clk(clk),
		.reset(rst),
		.din0(addsubIn3a),
		.din1(addsubIn3b),
		.opcode(addsubMod3),
		.ce(1'b1),
		.dout(addsubOut3Next)
	);
	reg [BitWidth-1:0] multIn0a, multIn0b;
	reg [BitWidth-1:0] multIn0aNext, multIn0bNext;
	wire [BitWidth-1:0] multOut0Next; reg [BitWidth-1:0] multOut0;
	iter_v2_fmul_32ns_32ns_32_10_full_dsp #(
		.ID(1),
		.NUM_STAGE(10),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_fmul_32ns_32ns_32_10_full_dsp_U0(
		.clk(clk),
		.reset(rst),
		.din0(multIn0a),
		.din1(multIn0b),
		.ce(1'b1),
		.dout(multOut0Next)
	);
	reg [BitWidth-1:0] multIn1a, multIn1b;
	reg [BitWidth-1:0] multIn1aNext, multIn1bNext;
	wire [BitWidth-1:0] multOut1Next; reg [BitWidth-1:0] multOut1;
	iter_v2_fmul_32ns_32ns_32_10_full_dsp #(
		.ID(1),
		.NUM_STAGE(10),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_fmul_32ns_32ns_32_10_full_dsp_U1(
		.clk(clk),
		.reset(rst),
		.din0(multIn1a),
		.din1(multIn1b),
		.ce(1'b1),
		.dout(multOut1Next)
	);
	reg [BitWidth-1:0] multIn2a, multIn2b;
	reg [BitWidth-1:0] multIn2aNext, multIn2bNext;
	wire [BitWidth-1:0] multOut2Next; reg [BitWidth-1:0] multOut2;
	iter_v2_fmul_32ns_32ns_32_10_full_dsp #(
		.ID(1),
		.NUM_STAGE(10),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_fmul_32ns_32ns_32_10_full_dsp_U2(
		.clk(clk),
		.reset(rst),
		.din0(multIn2a),
		.din1(multIn2b),
		.ce(1'b1),
		.dout(multOut2Next)
	);
	reg [BitWidth-1:0] divIn0a, divIn0b;
	reg [BitWidth-1:0] divIn0aNext, divIn0bNext;
	wire [BitWidth-1:0] divOut0Next; reg [BitWidth-1:0] divOut0;
	iter_v2_fdiv_32ns_32ns_32_30 #(
		.ID(1),
		.NUM_STAGE(30),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_fdiv_32ns_32ns_32_30_U0(
		.clk(clk),
		.reset(rst),
		.din0(divIn0a),
		.din1(divIn0b),
		.ce(1'b1),
		.dout(divOut0Next)
	);
	reg [BitWidth-1:0] sqrtIn0a;
	reg [BitWidth-1:0] sqrtIn0aNext;
	wire [BitWidth-1:0] sqrtOut0Next; reg [BitWidth-1:0] sqrtOut0;
	iter_v2_fsqrt_32ns_32ns_32_30 #(
		.ID(1),
		.NUM_STAGE(30),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(32))
	iter_v2_fsqrt_32ns_32ns_32_30_U0(
		.clk(clk),
		.reset(rst),
		.din0(0),
		.din1(sqrtIn0a),
		.ce(1'b1),
		.dout(sqrtOut0Next)
	);
	reg [BitWidth-1:0] eqgtgeltleneIn0a, eqgtgeltleneIn0b;
	reg [BitWidth-1:0] eqgtgeltleneMod0Next; reg [BitWidth-1:0] eqgtgeltleneMod0;
	reg [BitWidth-1:0] eqgtgeltleneIn0aNext, eqgtgeltleneIn0bNext;
	wire [BitWidth-1:0] eqgtgeltleneOut0Next; reg [BitWidth-1:0] eqgtgeltleneOut0;
	iter_v2_fcmp_32ns_32ns_1_4 #(
		.ID(1),
		.NUM_STAGE(4),
		.din0_WIDTH(32),
		.din1_WIDTH(32),
		.dout_WIDTH(1))
	iter_v2_fcmp_32ns_32ns_1_4_U0(
		.clk(clk),
		.reset(rst),
		.din0(eqgtgeltleneIn0a),
		.din1(eqgtgeltleneIn0b),
		.ce(1'b1),
		.opcode(eqgtgeltleneMod0),
		.dout(eqgtgeltleneOut0Next)
	);
	always@(posedge clk) begin
		addsubIn0a <= addsubIn0aNext;
		addsubIn0b <= addsubIn0bNext;
		addsubMod0 <= addsubMod0Next;
		addsubOut0 <= addsubOut0Next;
		addsubIn1a <= addsubIn1aNext;
		addsubIn1b <= addsubIn1bNext;
		addsubMod1 <= addsubMod1Next;
		addsubOut1 <= addsubOut1Next;
		addsubIn2a <= addsubIn2aNext;
		addsubIn2b <= addsubIn2bNext;
		addsubMod2 <= addsubMod2Next;
		addsubOut2 <= addsubOut2Next;
		addsubIn3a <= addsubIn3aNext;
		addsubIn3b <= addsubIn3bNext;
		addsubMod3 <= addsubMod3Next;
		addsubOut3 <= addsubOut3Next;
		multIn0a <= multIn0aNext;
		multIn0b <= multIn0bNext;
		multOut0 <= multOut0Next;
		multIn1a <= multIn1aNext;
		multIn1b <= multIn1bNext;
		multOut1 <= multOut1Next;
		multIn2a <= multIn2aNext;
		multIn2b <= multIn2bNext;
		multOut2 <= multOut2Next;
		divIn0a <= divIn0aNext;
		divIn0b <= divIn0bNext;
		divOut0 <= divOut0Next;
		sqrtIn0a <= sqrtIn0aNext;
		sqrtOut0 <= sqrtOut0Next;
		eqgtgeltleneIn0a <= eqgtgeltleneIn0aNext;
		eqgtgeltleneIn0b <= eqgtgeltleneIn0bNext;
		eqgtgeltleneMod0 <= eqgtgeltleneMod0Next;
		eqgtgeltleneOut0 <= eqgtgeltleneOut0Next;
		reg000 <= reg000Next; reg001 <= reg001Next; reg002 <= reg002Next; reg003 <= reg003Next; reg004 <= reg004Next; reg005 <= reg005Next; reg006 <= reg006Next; reg007 <= reg007Next; reg008 <= reg008Next; reg009 <= reg009Next; reg010 <= reg010Next; reg011 <= reg011Next; reg012 <= reg012Next; reg013 <= reg013Next; reg014 <= reg014Next; reg015 <= reg015Next; reg016 <= reg016Next; reg017 <= reg017Next; reg018 <= reg018Next; reg019 <= reg019Next; 
		reg020 <= reg020Next; reg021 <= reg021Next; reg022 <= reg022Next; reg023 <= reg023Next; reg024 <= reg024Next; reg025 <= reg025Next; reg026 <= reg026Next; reg027 <= reg027Next; reg028 <= reg028Next; reg029 <= reg029Next; reg030 <= reg030Next; reg031 <= reg031Next; reg032 <= reg032Next; reg033 <= reg033Next; reg034 <= reg034Next; reg035 <= reg035Next; reg036 <= reg036Next; reg037 <= reg037Next; reg038 <= reg038Next; reg039 <= reg039Next; 
		reg040 <= reg040Next; reg041 <= reg041Next; reg042 <= reg042Next; reg043 <= reg043Next; reg044 <= reg044Next; reg045 <= reg045Next; reg046 <= reg046Next; reg047 <= reg047Next; reg048 <= reg048Next; reg049 <= reg049Next; reg050 <= reg050Next; reg051 <= reg051Next; reg052 <= reg052Next; reg053 <= reg053Next; reg054 <= reg054Next; reg055 <= reg055Next; reg056 <= reg056Next; reg057 <= reg057Next; reg058 <= reg058Next; reg059 <= reg059Next; 
		reg060 <= reg060Next; reg061 <= reg061Next; reg062 <= reg062Next; reg063 <= reg063Next; reg064 <= reg064Next; reg065 <= reg065Next; reg066 <= reg066Next; reg067 <= reg067Next; reg068 <= reg068Next; reg069 <= reg069Next; reg070 <= reg070Next; reg071 <= reg071Next; reg072 <= reg072Next; reg073 <= reg073Next; reg074 <= reg074Next; reg075 <= reg075Next; reg076 <= reg076Next; reg077 <= reg077Next; reg078 <= reg078Next; reg079 <= reg079Next; 
		reg080 <= reg080Next; reg081 <= reg081Next; reg082 <= reg082Next; reg083 <= reg083Next; reg084 <= reg084Next; reg085 <= reg085Next; reg086 <= reg086Next; reg087 <= reg087Next; reg088 <= reg088Next; reg089 <= reg089Next; reg090 <= reg090Next; reg091 <= reg091Next; reg092 <= reg092Next; reg093 <= reg093Next; reg094 <= reg094Next; reg095 <= reg095Next; reg096 <= reg096Next; reg097 <= reg097Next; reg098 <= reg098Next; reg099 <= reg099Next; 
		reg100 <= reg100Next; reg101 <= reg101Next; reg102 <= reg102Next; reg103 <= reg103Next; reg104 <= reg104Next; reg105 <= reg105Next; reg106 <= reg106Next; reg107 <= reg107Next; reg108 <= reg108Next; reg109 <= reg109Next; reg110 <= reg110Next; reg111 <= reg111Next; reg112 <= reg112Next; reg113 <= reg113Next; reg114 <= reg114Next; reg115 <= reg115Next; reg116 <= reg116Next; reg117 <= reg117Next; reg118 <= reg118Next; reg119 <= reg119Next; 
		reg120 <= reg120Next; reg121 <= reg121Next; reg122 <= reg122Next; reg123 <= reg123Next; reg124 <= reg124Next; reg125 <= reg125Next; reg126 <= reg126Next; reg127 <= reg127Next; reg128 <= reg128Next; reg129 <= reg129Next; reg130 <= reg130Next; reg131 <= reg131Next; reg132 <= reg132Next; reg133 <= reg133Next; reg134 <= reg134Next; reg135 <= reg135Next; reg136 <= reg136Next; reg137 <= reg137Next; reg138 <= reg138Next; reg139 <= reg139Next; 
		reg140 <= reg140Next; reg141 <= reg141Next; reg142 <= reg142Next; reg143 <= reg143Next; reg144 <= reg144Next; reg145 <= reg145Next; reg146 <= reg146Next; reg147 <= reg147Next; reg148 <= reg148Next; reg149 <= reg149Next; reg150 <= reg150Next; reg151 <= reg151Next; reg152 <= reg152Next; reg153 <= reg153Next; reg154 <= reg154Next; reg155 <= reg155Next; reg156 <= reg156Next; reg157 <= reg157Next; reg158 <= reg158Next; reg159 <= reg159Next; 
		reg160 <= reg160Next; reg161 <= reg161Next; reg162 <= reg162Next; reg163 <= reg163Next; reg164 <= reg164Next; reg165 <= reg165Next; reg166 <= reg166Next; reg167 <= reg167Next; reg168 <= reg168Next; reg169 <= reg169Next; reg170 <= reg170Next; reg171 <= reg171Next; reg172 <= reg172Next; reg173 <= reg173Next; reg174 <= reg174Next; reg175 <= reg175Next; reg176 <= reg176Next; reg177 <= reg177Next; reg178 <= reg178Next; reg179 <= reg179Next; 
		reg180 <= reg180Next; reg181 <= reg181Next; reg182 <= reg182Next; reg183 <= reg183Next; reg184 <= reg184Next; reg185 <= reg185Next; reg186 <= reg186Next; reg187 <= reg187Next; reg188 <= reg188Next; reg189 <= reg189Next; reg190 <= reg190Next; reg191 <= reg191Next; reg192 <= reg192Next; reg193 <= reg193Next; reg194 <= reg194Next; reg195 <= reg195Next; reg196 <= reg196Next; reg197 <= reg197Next; reg198 <= reg198Next; reg199 <= reg199Next; 
		reg200 <= reg200Next; reg201 <= reg201Next; reg202 <= reg202Next; reg203 <= reg203Next; reg204 <= reg204Next; reg205 <= reg205Next; reg206 <= reg206Next; reg207 <= reg207Next; reg208 <= reg208Next; reg209 <= reg209Next; reg210 <= reg210Next; reg211 <= reg211Next; reg212 <= reg212Next; reg213 <= reg213Next; reg214 <= reg214Next; reg215 <= reg215Next; reg216 <= reg216Next; reg217 <= reg217Next; reg218 <= reg218Next; reg219 <= reg219Next; 
		reg220 <= reg220Next; reg221 <= reg221Next; reg222 <= reg222Next; reg223 <= reg223Next; reg224 <= reg224Next; reg225 <= reg225Next; reg226 <= reg226Next; reg227 <= reg227Next; reg228 <= reg228Next; reg229 <= reg229Next; reg230 <= reg230Next; reg231 <= reg231Next; reg232 <= reg232Next; reg233 <= reg233Next; reg234 <= reg234Next; reg235 <= reg235Next; reg236 <= reg236Next; reg237 <= reg237Next; reg238 <= reg238Next; reg239 <= reg239Next; 
		reg240 <= reg240Next; reg241 <= reg241Next; reg242 <= reg242Next; reg243 <= reg243Next; reg244 <= reg244Next; reg245 <= reg245Next; reg246 <= reg246Next; reg247 <= reg247Next; reg248 <= reg248Next; reg249 <= reg249Next; reg250 <= reg250Next; reg251 <= reg251Next; reg252 <= reg252Next; reg253 <= reg253Next; reg254 <= reg254Next; reg255 <= reg255Next; reg256 <= reg256Next; reg257 <= reg257Next; reg258 <= reg258Next; reg259 <= reg259Next; 
		reg260 <= reg260Next; reg261 <= reg261Next; reg262 <= reg262Next; reg263 <= reg263Next; reg264 <= reg264Next; reg265 <= reg265Next; reg266 <= reg266Next; reg267 <= reg267Next; reg268 <= reg268Next; reg269 <= reg269Next; reg270 <= reg270Next; reg271 <= reg271Next; reg272 <= reg272Next; reg273 <= reg273Next; reg274 <= reg274Next; reg275 <= reg275Next; reg276 <= reg276Next; reg277 <= reg277Next; reg278 <= reg278Next; reg279 <= reg279Next; 
		reg280 <= reg280Next; reg281 <= reg281Next; reg282 <= reg282Next; reg283 <= reg283Next; reg284 <= reg284Next; reg285 <= reg285Next; reg286 <= reg286Next; reg287 <= reg287Next; reg288 <= reg288Next; reg289 <= reg289Next; reg290 <= reg290Next; reg291 <= reg291Next; reg292 <= reg292Next; reg293 <= reg293Next; reg294 <= reg294Next; reg295 <= reg295Next; reg296 <= reg296Next; reg297 <= reg297Next; reg298 <= reg298Next; reg299 <= reg299Next; 
		reg300 <= reg300Next; reg301 <= reg301Next; reg302 <= reg302Next; reg303 <= reg303Next; reg304 <= reg304Next; reg305 <= reg305Next; reg306 <= reg306Next; reg307 <= reg307Next; reg308 <= reg308Next; reg309 <= reg309Next; reg310 <= reg310Next; reg311 <= reg311Next; reg312 <= reg312Next; reg313 <= reg313Next; reg314 <= reg314Next; reg315 <= reg315Next; reg316 <= reg316Next; reg317 <= reg317Next; reg318 <= reg318Next; reg319 <= reg319Next; 
		reg320 <= reg320Next; reg321 <= reg321Next; reg322 <= reg322Next; reg323 <= reg323Next; reg324 <= reg324Next; reg325 <= reg325Next; reg326 <= reg326Next; reg327 <= reg327Next; reg328 <= reg328Next; reg329 <= reg329Next; reg330 <= reg330Next; reg331 <= reg331Next; reg332 <= reg332Next; reg333 <= reg333Next; reg334 <= reg334Next; reg335 <= reg335Next; reg336 <= reg336Next; reg337 <= reg337Next; reg338 <= reg338Next; reg339 <= reg339Next; 
		reg340 <= reg340Next; reg341 <= reg341Next; reg342 <= reg342Next; reg343 <= reg343Next; reg344 <= reg344Next; reg345 <= reg345Next; reg346 <= reg346Next; reg347 <= reg347Next; reg348 <= reg348Next; reg349 <= reg349Next; reg350 <= reg350Next; reg351 <= reg351Next; reg352 <= reg352Next; reg353 <= reg353Next; reg354 <= reg354Next; reg355 <= reg355Next; reg356 <= reg356Next; reg357 <= reg357Next; reg358 <= reg358Next; reg359 <= reg359Next; 
		reg360 <= reg360Next; reg361 <= reg361Next; reg362 <= reg362Next; reg363 <= reg363Next; reg364 <= reg364Next; reg365 <= reg365Next; reg366 <= reg366Next; reg367 <= reg367Next; reg368 <= reg368Next; reg369 <= reg369Next; reg370 <= reg370Next; reg371 <= reg371Next; reg372 <= reg372Next; reg373 <= reg373Next; reg374 <= reg374Next; reg375 <= reg375Next; reg376 <= reg376Next; reg377 <= reg377Next; reg378 <= reg378Next; reg379 <= reg379Next; 
		reg380 <= reg380Next; reg381 <= reg381Next; reg382 <= reg382Next; reg383 <= reg383Next; reg384 <= reg384Next; reg385 <= reg385Next; reg386 <= reg386Next; reg387 <= reg387Next; reg388 <= reg388Next; reg389 <= reg389Next; reg390 <= reg390Next; reg391 <= reg391Next; reg392 <= reg392Next; reg393 <= reg393Next; reg394 <= reg394Next; reg395 <= reg395Next; reg396 <= reg396Next; reg397 <= reg397Next; reg398 <= reg398Next; reg399 <= reg399Next; 
		reg400 <= reg400Next; reg401 <= reg401Next; reg402 <= reg402Next; reg403 <= reg403Next; reg404 <= reg404Next; reg405 <= reg405Next; reg406 <= reg406Next; reg407 <= reg407Next; reg408 <= reg408Next; reg409 <= reg409Next; reg410 <= reg410Next; reg411 <= reg411Next; reg412 <= reg412Next; reg413 <= reg413Next; reg414 <= reg414Next; reg415 <= reg415Next; reg416 <= reg416Next; reg417 <= reg417Next; reg418 <= reg418Next; reg419 <= reg419Next; 
		reg420 <= reg420Next; reg421 <= reg421Next; reg422 <= reg422Next; reg423 <= reg423Next; reg424 <= reg424Next; reg425 <= reg425Next; reg426 <= reg426Next; reg427 <= reg427Next; reg428 <= reg428Next; reg429 <= reg429Next; reg430 <= reg430Next; reg431 <= reg431Next; reg432 <= reg432Next; reg433 <= reg433Next; reg434 <= reg434Next; reg435 <= reg435Next; reg436 <= reg436Next; reg437 <= reg437Next; reg438 <= reg438Next; reg439 <= reg439Next; 
		reg440 <= reg440Next; reg441 <= reg441Next; reg442 <= reg442Next; reg443 <= reg443Next; reg444 <= reg444Next; reg445 <= reg445Next; reg446 <= reg446Next; reg447 <= reg447Next; reg448 <= reg448Next; reg449 <= reg449Next; reg450 <= reg450Next; reg451 <= reg451Next; reg452 <= reg452Next; reg453 <= reg453Next; reg454 <= reg454Next; reg455 <= reg455Next; reg456 <= reg456Next; reg457 <= reg457Next; reg458 <= reg458Next; reg459 <= reg459Next; 
		reg460 <= reg460Next; reg461 <= reg461Next; reg462 <= reg462Next; reg463 <= reg463Next; reg464 <= reg464Next; reg465 <= reg465Next; reg466 <= reg466Next; reg467 <= reg467Next; reg468 <= reg468Next; reg469 <= reg469Next; reg470 <= reg470Next; reg471 <= reg471Next; reg472 <= reg472Next; reg473 <= reg473Next; reg474 <= reg474Next; reg475 <= reg475Next; reg476 <= reg476Next; reg477 <= reg477Next; reg478 <= reg478Next; reg479 <= reg479Next; 
		reg480 <= reg480Next; reg481 <= reg481Next; reg482 <= reg482Next; reg483 <= reg483Next; reg484 <= reg484Next; reg485 <= reg485Next; reg486 <= reg486Next; reg487 <= reg487Next; reg488 <= reg488Next; reg489 <= reg489Next; reg490 <= reg490Next; reg491 <= reg491Next; reg492 <= reg492Next; reg493 <= reg493Next; reg494 <= reg494Next; reg495 <= reg495Next; reg496 <= reg496Next; reg497 <= reg497Next; reg498 <= reg498Next; reg499 <= reg499Next; 
		reg500 <= reg500Next; reg501 <= reg501Next; reg502 <= reg502Next; reg503 <= reg503Next; reg504 <= reg504Next; reg505 <= reg505Next; reg506 <= reg506Next; reg507 <= reg507Next; reg508 <= reg508Next; reg509 <= reg509Next; reg510 <= reg510Next; reg511 <= reg511Next; reg512 <= reg512Next; reg513 <= reg513Next; reg514 <= reg514Next; reg515 <= reg515Next; reg516 <= reg516Next; reg517 <= reg517Next; reg518 <= reg518Next; reg519 <= reg519Next; 
		reg520 <= reg520Next; reg521 <= reg521Next; reg522 <= reg522Next; reg523 <= reg523Next; reg524 <= reg524Next; reg525 <= reg525Next; reg526 <= reg526Next; reg527 <= reg527Next; reg528 <= reg528Next; reg529 <= reg529Next; reg530 <= reg530Next; reg531 <= reg531Next; reg532 <= reg532Next; reg533 <= reg533Next; reg534 <= reg534Next; reg535 <= reg535Next; reg536 <= reg536Next; reg537 <= reg537Next; reg538 <= reg538Next; reg539 <= reg539Next; 
		reg540 <= reg540Next; reg541 <= reg541Next; reg542 <= reg542Next; reg543 <= reg543Next; reg544 <= reg544Next; reg545 <= reg545Next; reg546 <= reg546Next; reg547 <= reg547Next; reg548 <= reg548Next; reg549 <= reg549Next; reg550 <= reg550Next; reg551 <= reg551Next; reg552 <= reg552Next; reg553 <= reg553Next; reg554 <= reg554Next; reg555 <= reg555Next; reg556 <= reg556Next; reg557 <= reg557Next; reg558 <= reg558Next; reg559 <= reg559Next; 
		reg560 <= reg560Next; reg561 <= reg561Next; reg562 <= reg562Next; reg563 <= reg563Next; reg564 <= reg564Next; reg565 <= reg565Next; reg566 <= reg566Next; reg567 <= reg567Next; reg568 <= reg568Next; reg569 <= reg569Next; reg570 <= reg570Next; reg571 <= reg571Next; reg572 <= reg572Next; reg573 <= reg573Next; reg574 <= reg574Next; reg575 <= reg575Next; reg576 <= reg576Next; reg577 <= reg577Next; reg578 <= reg578Next; reg579 <= reg579Next; 
		reg580 <= reg580Next; reg581 <= reg581Next; reg582 <= reg582Next; reg583 <= reg583Next; reg584 <= reg584Next; reg585 <= reg585Next; reg586 <= reg586Next; reg587 <= reg587Next; reg588 <= reg588Next; reg589 <= reg589Next; reg590 <= reg590Next; reg591 <= reg591Next; reg592 <= reg592Next; reg593 <= reg593Next; reg594 <= reg594Next; reg595 <= reg595Next; reg596 <= reg596Next; reg597 <= reg597Next; reg598 <= reg598Next; reg599 <= reg599Next; 
		reg600 <= reg600Next; reg601 <= reg601Next; reg602 <= reg602Next; reg603 <= reg603Next; reg604 <= reg604Next; reg605 <= reg605Next; reg606 <= reg606Next; reg607 <= reg607Next; reg608 <= reg608Next; reg609 <= reg609Next; reg610 <= reg610Next; reg611 <= reg611Next; reg612 <= reg612Next; reg613 <= reg613Next; reg614 <= reg614Next; reg615 <= reg615Next; reg616 <= reg616Next; reg617 <= reg617Next; reg618 <= reg618Next; reg619 <= reg619Next; 
		reg620 <= reg620Next; reg621 <= reg621Next; reg622 <= reg622Next; reg623 <= reg623Next; reg624 <= reg624Next; reg625 <= reg625Next; reg626 <= reg626Next; reg627 <= reg627Next; reg628 <= reg628Next; reg629 <= reg629Next; reg630 <= reg630Next; reg631 <= reg631Next; reg632 <= reg632Next; reg633 <= reg633Next; reg634 <= reg634Next; reg635 <= reg635Next; reg636 <= reg636Next; reg637 <= reg637Next; reg638 <= reg638Next; reg639 <= reg639Next; 
		reg640 <= reg640Next; reg641 <= reg641Next; reg642 <= reg642Next; reg643 <= reg643Next; reg644 <= reg644Next; reg645 <= reg645Next; reg646 <= reg646Next; reg647 <= reg647Next; reg648 <= reg648Next; reg649 <= reg649Next; reg650 <= reg650Next; reg651 <= reg651Next; reg652 <= reg652Next; reg653 <= reg653Next; reg654 <= reg654Next; reg655 <= reg655Next; reg656 <= reg656Next; reg657 <= reg657Next; reg658 <= reg658Next; reg659 <= reg659Next; 
		reg660 <= reg660Next; reg661 <= reg661Next; reg662 <= reg662Next; reg663 <= reg663Next; reg664 <= reg664Next; reg665 <= reg665Next; reg666 <= reg666Next; reg667 <= reg667Next; reg668 <= reg668Next; reg669 <= reg669Next; reg670 <= reg670Next; reg671 <= reg671Next; reg672 <= reg672Next; reg673 <= reg673Next; reg674 <= reg674Next; reg675 <= reg675Next; reg676 <= reg676Next; reg677 <= reg677Next; reg678 <= reg678Next; reg679 <= reg679Next; 
		reg680 <= reg680Next; reg681 <= reg681Next; reg682 <= reg682Next; reg683 <= reg683Next; reg684 <= reg684Next; reg685 <= reg685Next; reg686 <= reg686Next; reg687 <= reg687Next; reg688 <= reg688Next; reg689 <= reg689Next; reg690 <= reg690Next; reg691 <= reg691Next; reg692 <= reg692Next; reg693 <= reg693Next; reg694 <= reg694Next; reg695 <= reg695Next; reg696 <= reg696Next; reg697 <= reg697Next; reg698 <= reg698Next; reg699 <= reg699Next; 
		reg700 <= reg700Next; reg701 <= reg701Next; reg702 <= reg702Next; reg703 <= reg703Next; reg704 <= reg704Next; reg705 <= reg705Next; reg706 <= reg706Next; reg707 <= reg707Next; reg708 <= reg708Next; reg709 <= reg709Next; reg710 <= reg710Next; reg711 <= reg711Next; reg712 <= reg712Next; reg713 <= reg713Next; reg714 <= reg714Next; reg715 <= reg715Next; reg716 <= reg716Next; reg717 <= reg717Next; reg718 <= reg718Next; 
	end
	always@(*) begin
		reg000Next = reg000; reg001Next = reg001; reg002Next = reg002; reg003Next = reg003; reg004Next = reg004; reg005Next = reg005; reg006Next = reg006; reg007Next = reg007; reg008Next = reg008; reg009Next = reg009; reg010Next = reg010; reg011Next = reg011; reg012Next = reg012; reg013Next = reg013; reg014Next = reg014; reg015Next = reg015; reg016Next = reg016; reg017Next = reg017; reg018Next = reg018; reg019Next = reg019; 
		reg020Next = reg020; reg021Next = reg021; reg022Next = reg022; reg023Next = reg023; reg024Next = reg024; reg025Next = reg025; reg026Next = reg026; reg027Next = reg027; reg028Next = reg028; reg029Next = reg029; reg030Next = reg030; reg031Next = reg031; reg032Next = reg032; reg033Next = reg033; reg034Next = reg034; reg035Next = reg035; reg036Next = reg036; reg037Next = reg037; reg038Next = reg038; reg039Next = reg039; 
		reg040Next = reg040; reg041Next = reg041; reg042Next = reg042; reg043Next = reg043; reg044Next = reg044; reg045Next = reg045; reg046Next = reg046; reg047Next = reg047; reg048Next = reg048; reg049Next = reg049; reg050Next = reg050; reg051Next = reg051; reg052Next = reg052; reg053Next = reg053; reg054Next = reg054; reg055Next = reg055; reg056Next = reg056; reg057Next = reg057; reg058Next = reg058; reg059Next = reg059; 
		reg060Next = reg060; reg061Next = reg061; reg062Next = reg062; reg063Next = reg063; reg064Next = reg064; reg065Next = reg065; reg066Next = reg066; reg067Next = reg067; reg068Next = reg068; reg069Next = reg069; reg070Next = reg070; reg071Next = reg071; reg072Next = reg072; reg073Next = reg073; reg074Next = reg074; reg075Next = reg075; reg076Next = reg076; reg077Next = reg077; reg078Next = reg078; reg079Next = reg079; 
		reg080Next = reg080; reg081Next = reg081; reg082Next = reg082; reg083Next = reg083; reg084Next = reg084; reg085Next = reg085; reg086Next = reg086; reg087Next = reg087; reg088Next = reg088; reg089Next = reg089; reg090Next = reg090; reg091Next = reg091; reg092Next = reg092; reg093Next = reg093; reg094Next = reg094; reg095Next = reg095; reg096Next = reg096; reg097Next = reg097; reg098Next = reg098; reg099Next = reg099; 
		reg100Next = reg100; reg101Next = reg101; reg102Next = reg102; reg103Next = reg103; reg104Next = reg104; reg105Next = reg105; reg106Next = reg106; reg107Next = reg107; reg108Next = reg108; reg109Next = reg109; reg110Next = reg110; reg111Next = reg111; reg112Next = reg112; reg113Next = reg113; reg114Next = reg114; reg115Next = reg115; reg116Next = reg116; reg117Next = reg117; reg118Next = reg118; reg119Next = reg119; 
		reg120Next = reg120; reg121Next = reg121; reg122Next = reg122; reg123Next = reg123; reg124Next = reg124; reg125Next = reg125; reg126Next = reg126; reg127Next = reg127; reg128Next = reg128; reg129Next = reg129; reg130Next = reg130; reg131Next = reg131; reg132Next = reg132; reg133Next = reg133; reg134Next = reg134; reg135Next = reg135; reg136Next = reg136; reg137Next = reg137; reg138Next = reg138; reg139Next = reg139; 
		reg140Next = reg140; reg141Next = reg141; reg142Next = reg142; reg143Next = reg143; reg144Next = reg144; reg145Next = reg145; reg146Next = reg146; reg147Next = reg147; reg148Next = reg148; reg149Next = reg149; reg150Next = reg150; reg151Next = reg151; reg152Next = reg152; reg153Next = reg153; reg154Next = reg154; reg155Next = reg155; reg156Next = reg156; reg157Next = reg157; reg158Next = reg158; reg159Next = reg159; 
		reg160Next = reg160; reg161Next = reg161; reg162Next = reg162; reg163Next = reg163; reg164Next = reg164; reg165Next = reg165; reg166Next = reg166; reg167Next = reg167; reg168Next = reg168; reg169Next = reg169; reg170Next = reg170; reg171Next = reg171; reg172Next = reg172; reg173Next = reg173; reg174Next = reg174; reg175Next = reg175; reg176Next = reg176; reg177Next = reg177; reg178Next = reg178; reg179Next = reg179; 
		reg180Next = reg180; reg181Next = reg181; reg182Next = reg182; reg183Next = reg183; reg184Next = reg184; reg185Next = reg185; reg186Next = reg186; reg187Next = reg187; reg188Next = reg188; reg189Next = reg189; reg190Next = reg190; reg191Next = reg191; reg192Next = reg192; reg193Next = reg193; reg194Next = reg194; reg195Next = reg195; reg196Next = reg196; reg197Next = reg197; reg198Next = reg198; reg199Next = reg199; 
		reg200Next = reg200; reg201Next = reg201; reg202Next = reg202; reg203Next = reg203; reg204Next = reg204; reg205Next = reg205; reg206Next = reg206; reg207Next = reg207; reg208Next = reg208; reg209Next = reg209; reg210Next = reg210; reg211Next = reg211; reg212Next = reg212; reg213Next = reg213; reg214Next = reg214; reg215Next = reg215; reg216Next = reg216; reg217Next = reg217; reg218Next = reg218; reg219Next = reg219; 
		reg220Next = reg220; reg221Next = reg221; reg222Next = reg222; reg223Next = reg223; reg224Next = reg224; reg225Next = reg225; reg226Next = reg226; reg227Next = reg227; reg228Next = reg228; reg229Next = reg229; reg230Next = reg230; reg231Next = reg231; reg232Next = reg232; reg233Next = reg233; reg234Next = reg234; reg235Next = reg235; reg236Next = reg236; reg237Next = reg237; reg238Next = reg238; reg239Next = reg239; 
		reg240Next = reg240; reg241Next = reg241; reg242Next = reg242; reg243Next = reg243; reg244Next = reg244; reg245Next = reg245; reg246Next = reg246; reg247Next = reg247; reg248Next = reg248; reg249Next = reg249; reg250Next = reg250; reg251Next = reg251; reg252Next = reg252; reg253Next = reg253; reg254Next = reg254; reg255Next = reg255; reg256Next = reg256; reg257Next = reg257; reg258Next = reg258; reg259Next = reg259; 
		reg260Next = reg260; reg261Next = reg261; reg262Next = reg262; reg263Next = reg263; reg264Next = reg264; reg265Next = reg265; reg266Next = reg266; reg267Next = reg267; reg268Next = reg268; reg269Next = reg269; reg270Next = reg270; reg271Next = reg271; reg272Next = reg272; reg273Next = reg273; reg274Next = reg274; reg275Next = reg275; reg276Next = reg276; reg277Next = reg277; reg278Next = reg278; reg279Next = reg279; 
		reg280Next = reg280; reg281Next = reg281; reg282Next = reg282; reg283Next = reg283; reg284Next = reg284; reg285Next = reg285; reg286Next = reg286; reg287Next = reg287; reg288Next = reg288; reg289Next = reg289; reg290Next = reg290; reg291Next = reg291; reg292Next = reg292; reg293Next = reg293; reg294Next = reg294; reg295Next = reg295; reg296Next = reg296; reg297Next = reg297; reg298Next = reg298; reg299Next = reg299; 
		reg300Next = reg300; reg301Next = reg301; reg302Next = reg302; reg303Next = reg303; reg304Next = reg304; reg305Next = reg305; reg306Next = reg306; reg307Next = reg307; reg308Next = reg308; reg309Next = reg309; reg310Next = reg310; reg311Next = reg311; reg312Next = reg312; reg313Next = reg313; reg314Next = reg314; reg315Next = reg315; reg316Next = reg316; reg317Next = reg317; reg318Next = reg318; reg319Next = reg319; 
		reg320Next = reg320; reg321Next = reg321; reg322Next = reg322; reg323Next = reg323; reg324Next = reg324; reg325Next = reg325; reg326Next = reg326; reg327Next = reg327; reg328Next = reg328; reg329Next = reg329; reg330Next = reg330; reg331Next = reg331; reg332Next = reg332; reg333Next = reg333; reg334Next = reg334; reg335Next = reg335; reg336Next = reg336; reg337Next = reg337; reg338Next = reg338; reg339Next = reg339; 
		reg340Next = reg340; reg341Next = reg341; reg342Next = reg342; reg343Next = reg343; reg344Next = reg344; reg345Next = reg345; reg346Next = reg346; reg347Next = reg347; reg348Next = reg348; reg349Next = reg349; reg350Next = reg350; reg351Next = reg351; reg352Next = reg352; reg353Next = reg353; reg354Next = reg354; reg355Next = reg355; reg356Next = reg356; reg357Next = reg357; reg358Next = reg358; reg359Next = reg359; 
		reg360Next = reg360; reg361Next = reg361; reg362Next = reg362; reg363Next = reg363; reg364Next = reg364; reg365Next = reg365; reg366Next = reg366; reg367Next = reg367; reg368Next = reg368; reg369Next = reg369; reg370Next = reg370; reg371Next = reg371; reg372Next = reg372; reg373Next = reg373; reg374Next = reg374; reg375Next = reg375; reg376Next = reg376; reg377Next = reg377; reg378Next = reg378; reg379Next = reg379; 
		reg380Next = reg380; reg381Next = reg381; reg382Next = reg382; reg383Next = reg383; reg384Next = reg384; reg385Next = reg385; reg386Next = reg386; reg387Next = reg387; reg388Next = reg388; reg389Next = reg389; reg390Next = reg390; reg391Next = reg391; reg392Next = reg392; reg393Next = reg393; reg394Next = reg394; reg395Next = reg395; reg396Next = reg396; reg397Next = reg397; reg398Next = reg398; reg399Next = reg399; 
		reg400Next = reg400; reg401Next = reg401; reg402Next = reg402; reg403Next = reg403; reg404Next = reg404; reg405Next = reg405; reg406Next = reg406; reg407Next = reg407; reg408Next = reg408; reg409Next = reg409; reg410Next = reg410; reg411Next = reg411; reg412Next = reg412; reg413Next = reg413; reg414Next = reg414; reg415Next = reg415; reg416Next = reg416; reg417Next = reg417; reg418Next = reg418; reg419Next = reg419; 
		reg420Next = reg420; reg421Next = reg421; reg422Next = reg422; reg423Next = reg423; reg424Next = reg424; reg425Next = reg425; reg426Next = reg426; reg427Next = reg427; reg428Next = reg428; reg429Next = reg429; reg430Next = reg430; reg431Next = reg431; reg432Next = reg432; reg433Next = reg433; reg434Next = reg434; reg435Next = reg435; reg436Next = reg436; reg437Next = reg437; reg438Next = reg438; reg439Next = reg439; 
		reg440Next = reg440; reg441Next = reg441; reg442Next = reg442; reg443Next = reg443; reg444Next = reg444; reg445Next = reg445; reg446Next = reg446; reg447Next = reg447; reg448Next = reg448; reg449Next = reg449; reg450Next = reg450; reg451Next = reg451; reg452Next = reg452; reg453Next = reg453; reg454Next = reg454; reg455Next = reg455; reg456Next = reg456; reg457Next = reg457; reg458Next = reg458; reg459Next = reg459; 
		reg460Next = reg460; reg461Next = reg461; reg462Next = reg462; reg463Next = reg463; reg464Next = reg464; reg465Next = reg465; reg466Next = reg466; reg467Next = reg467; reg468Next = reg468; reg469Next = reg469; reg470Next = reg470; reg471Next = reg471; reg472Next = reg472; reg473Next = reg473; reg474Next = reg474; reg475Next = reg475; reg476Next = reg476; reg477Next = reg477; reg478Next = reg478; reg479Next = reg479; 
		reg480Next = reg480; reg481Next = reg481; reg482Next = reg482; reg483Next = reg483; reg484Next = reg484; reg485Next = reg485; reg486Next = reg486; reg487Next = reg487; reg488Next = reg488; reg489Next = reg489; reg490Next = reg490; reg491Next = reg491; reg492Next = reg492; reg493Next = reg493; reg494Next = reg494; reg495Next = reg495; reg496Next = reg496; reg497Next = reg497; reg498Next = reg498; reg499Next = reg499; 
		reg500Next = reg500; reg501Next = reg501; reg502Next = reg502; reg503Next = reg503; reg504Next = reg504; reg505Next = reg505; reg506Next = reg506; reg507Next = reg507; reg508Next = reg508; reg509Next = reg509; reg510Next = reg510; reg511Next = reg511; reg512Next = reg512; reg513Next = reg513; reg514Next = reg514; reg515Next = reg515; reg516Next = reg516; reg517Next = reg517; reg518Next = reg518; reg519Next = reg519; 
		reg520Next = reg520; reg521Next = reg521; reg522Next = reg522; reg523Next = reg523; reg524Next = reg524; reg525Next = reg525; reg526Next = reg526; reg527Next = reg527; reg528Next = reg528; reg529Next = reg529; reg530Next = reg530; reg531Next = reg531; reg532Next = reg532; reg533Next = reg533; reg534Next = reg534; reg535Next = reg535; reg536Next = reg536; reg537Next = reg537; reg538Next = reg538; reg539Next = reg539; 
		reg540Next = reg540; reg541Next = reg541; reg542Next = reg542; reg543Next = reg543; reg544Next = reg544; reg545Next = reg545; reg546Next = reg546; reg547Next = reg547; reg548Next = reg548; reg549Next = reg549; reg550Next = reg550; reg551Next = reg551; reg552Next = reg552; reg553Next = reg553; reg554Next = reg554; reg555Next = reg555; reg556Next = reg556; reg557Next = reg557; reg558Next = reg558; reg559Next = reg559; 
		reg560Next = reg560; reg561Next = reg561; reg562Next = reg562; reg563Next = reg563; reg564Next = reg564; reg565Next = reg565; reg566Next = reg566; reg567Next = reg567; reg568Next = reg568; reg569Next = reg569; reg570Next = reg570; reg571Next = reg571; reg572Next = reg572; reg573Next = reg573; reg574Next = reg574; reg575Next = reg575; reg576Next = reg576; reg577Next = reg577; reg578Next = reg578; reg579Next = reg579; 
		reg580Next = reg580; reg581Next = reg581; reg582Next = reg582; reg583Next = reg583; reg584Next = reg584; reg585Next = reg585; reg586Next = reg586; reg587Next = reg587; reg588Next = reg588; reg589Next = reg589; reg590Next = reg590; reg591Next = reg591; reg592Next = reg592; reg593Next = reg593; reg594Next = reg594; reg595Next = reg595; reg596Next = reg596; reg597Next = reg597; reg598Next = reg598; reg599Next = reg599; 
		reg600Next = reg600; reg601Next = reg601; reg602Next = reg602; reg603Next = reg603; reg604Next = reg604; reg605Next = reg605; reg606Next = reg606; reg607Next = reg607; reg608Next = reg608; reg609Next = reg609; reg610Next = reg610; reg611Next = reg611; reg612Next = reg612; reg613Next = reg613; reg614Next = reg614; reg615Next = reg615; reg616Next = reg616; reg617Next = reg617; reg618Next = reg618; reg619Next = reg619; 
		reg620Next = reg620; reg621Next = reg621; reg622Next = reg622; reg623Next = reg623; reg624Next = reg624; reg625Next = reg625; reg626Next = reg626; reg627Next = reg627; reg628Next = reg628; reg629Next = reg629; reg630Next = reg630; reg631Next = reg631; reg632Next = reg632; reg633Next = reg633; reg634Next = reg634; reg635Next = reg635; reg636Next = reg636; reg637Next = reg637; reg638Next = reg638; reg639Next = reg639; 
		reg640Next = reg640; reg641Next = reg641; reg642Next = reg642; reg643Next = reg643; reg644Next = reg644; reg645Next = reg645; reg646Next = reg646; reg647Next = reg647; reg648Next = reg648; reg649Next = reg649; reg650Next = reg650; reg651Next = reg651; reg652Next = reg652; reg653Next = reg653; reg654Next = reg654; reg655Next = reg655; reg656Next = reg656; reg657Next = reg657; reg658Next = reg658; reg659Next = reg659; 
		reg660Next = reg660; reg661Next = reg661; reg662Next = reg662; reg663Next = reg663; reg664Next = reg664; reg665Next = reg665; reg666Next = reg666; reg667Next = reg667; reg668Next = reg668; reg669Next = reg669; reg670Next = reg670; reg671Next = reg671; reg672Next = reg672; reg673Next = reg673; reg674Next = reg674; reg675Next = reg675; reg676Next = reg676; reg677Next = reg677; reg678Next = reg678; reg679Next = reg679; 
		reg680Next = reg680; reg681Next = reg681; reg682Next = reg682; reg683Next = reg683; reg684Next = reg684; reg685Next = reg685; reg686Next = reg686; reg687Next = reg687; reg688Next = reg688; reg689Next = reg689; reg690Next = reg690; reg691Next = reg691; reg692Next = reg692; reg693Next = reg693; reg694Next = reg694; reg695Next = reg695; reg696Next = reg696; reg697Next = reg697; reg698Next = reg698; reg699Next = reg699; 
		reg700Next = reg700; reg701Next = reg701; reg702Next = reg702; reg703Next = reg703; reg704Next = reg704; reg705Next = reg705; reg706Next = reg706; reg707Next = reg707; reg708Next = reg708; reg709Next = reg709; reg710Next = reg710; reg711Next = reg711; reg712Next = reg712; reg713Next = reg713; reg714Next = reg714; reg715Next = reg715; reg716Next = reg716; reg717Next = reg717; reg718Next = reg718; 
		addsubIn0aNext = 'bx;
		addsubIn0bNext = 'bx;
		addsubMod0Next = 'bx;
		addsubIn1aNext = 'bx;
		addsubIn1bNext = 'bx;
		addsubMod1Next = 'bx;
		addsubIn2aNext = 'bx;
		addsubIn2bNext = 'bx;
		addsubMod2Next = 'bx;
		addsubIn3aNext = 'bx;
		addsubIn3bNext = 'bx;
		addsubMod3Next = 'bx;
		multIn0aNext = 'bx;
		multIn0bNext = 'bx;
		multIn1aNext = 'bx;
		multIn1bNext = 'bx;
		multIn2aNext = 'bx;
		multIn2bNext = 'bx;
		divIn0aNext = 'bx;
		divIn0bNext = 'bx;
		sqrtIn0aNext = 'bx;
		eqgtgeltleneIn0aNext = 'bx;
		eqgtgeltleneIn0bNext = 'bx;
		eqgtgeltleneMod0Next = 'bx;
		uOut = addsubOut1;
		u_Out = addsubOut1;
		vOut = addsubOut2;
		v_Out = addsubOut2;
		wOut = addsubOut3;
		w_Out = addsubOut3;
		p3Out = divOut0;
		p4Out = divOut0;
		p5Out = divOut0;
		p0Out = divOut0;
		p2Out = divOut0;
		p1Out = divOut0;
		case(state)
		0:begin
			// s000
			addsubIn0aNext = u_S1; addsubIn0bNext = u_S0; addsubMod0Next = sub; 
			// s100
			addsubIn1aNext = v_S1; addsubIn1bNext = v_S0; addsubMod1Next = sub; 
			// s200
			addsubIn2aNext = w_S1; addsubIn2bNext = w_S0; addsubMod2Next = sub; 
			// s300
			addsubIn3aNext = u_S2; addsubIn3bNext = u_S0; addsubMod3Next = sub; 
			// cons1
			multIn0aNext = cons0; multIn0bNext = I_grad_sqrS; 
			// cons3
			multIn1aNext = cons0; multIn1bNext = I_xS; 
			// cons4
			multIn2aNext = cons0; multIn2bNext = I_yS; 
			// d074
			divIn0aNext = reg434; divIn0bNext = reg449; 
			// c080
			eqgtgeltleneIn0aNext = addsubOut3; eqgtgeltleneIn0bNext = reg559; eqgtgeltleneMod0Next = lt; 
			// d041
			reg450Next = divOut0;
			// s223
			reg454Next = addsubOut0;
			// m035
			reg456Next = multOut0;
			// m046
			reg457Next = multOut1;
			// m202
			reg490Next = multOut2;
			// a158
			reg494Next = addsubOut1;
			// a257
			reg495Next = addsubOut2;
			// a374
			reg500Next = addsubOut3;
			reg000Next = v_S0;
			reg001Next = w_S0;
			reg002Next = p0;
			reg005Next = p2;
			reg008Next = p4;
			reg011Next = jj;
			reg033Next = v_S2;
			reg034Next = w_S2;
			reg035Next = p1;
			reg038Next = p3;
			reg041Next = p5;
			reg044Next = ii;
			reg066Next = p0Prev;
			reg082Next = p2Prev;
			reg099Next = p4Prev;
			reg114Next = p1S_1;
			reg131Next = p3S_1;
			reg148Next = p5S_1;
			reg163Next = uS;
			reg198Next = vS;
			reg233Next = wS;
			reg268Next = u0S;
			reg291Next = v0S;
			reg315Next = I_xS;
			reg339Next = I_yS;
			reg364Next = I_tS;
			reg387Next = I_grad_sqrS;
			reg388Next = beta;
		end
		1:begin
			// s400
			addsubIn0aNext = reg033; addsubIn0bNext = reg000; addsubMod0Next = sub; 
			// s011
			addsubIn1aNext = reg034; addsubIn1bNext = reg001; addsubMod1Next = sub; 
			// s096
			addsubIn2aNext = reg098; addsubIn2bNext = reg450; addsubMod2Next = sub; 
			if ( reg060 != 0 && reg027 == 0 ) begin
				addsubIn2aNext = ZERO; addsubIn2bNext = reg450; addsubMod2Next = sub; 
			end
			// s087
			addsubIn3aNext = reg130; addsubIn3bNext = divOut0; addsubMod3Next = sub; 
			if ( reg060 == 0 && reg027 != 0 ) begin
				addsubIn3aNext = ZERO; addsubIn3bNext = divOut0; addsubMod3Next = sub; 
			end
			// m283
			multIn0aNext = reg500; multIn0bNext = reg591; 
			// m382
			multIn1aNext = reg500; multIn1bNext = reg619; 
			// m482
			multIn2aNext = reg500; multIn2bNext = reg647; 
			// d052
			divIn0aNext = reg414; divIn0bNext = sqrtOut0; 
			// c091
			eqgtgeltleneIn0aNext = reg500; eqgtgeltleneIn0bNext = reg530; eqgtgeltleneMod0Next = gt; 
			// ct0
			reg447Next = sqrtOut0;
			// s058
			reg458Next = addsubOut0;
			// m182
			reg491Next = multOut0;
			// m103
			reg493Next = multOut1;
			// as335
			reg713Next = addsubOut1;
			// as432
			reg714Next = addsubOut2;
			// as049
			reg715Next = addsubOut3;
		end
		2:begin
			// s212
			addsubIn0aNext = reg147; addsubIn0bNext = divOut0; addsubMod0Next = sub; 
			if ( reg060 == 0 && reg027 != 0 ) begin
				addsubIn0aNext = ZERO; addsubIn0bNext = divOut0; addsubMod0Next = sub; 
			end
			// a234
			addsubIn1aNext = reg453; addsubIn1bNext = reg454; addsubMod1Next = add; 
			// s187
			addsubIn2aNext = reg219; addsubIn2bNext = reg456; addsubMod2Next = sub; 
			if ( reg065 == 0 && reg032 == 0 ) begin
				addsubIn2aNext = reg219; addsubIn2bNext = ZERO; addsubMod2Next = sub; 
			end
			// s295
			addsubIn3aNext = reg252; addsubIn3bNext = reg457; addsubMod3Next = sub; 
			if ( reg063 == 0 && reg030 == 0 ) begin
				addsubIn3aNext = reg252; addsubIn3bNext = ZERO; addsubMod3Next = sub; 
			end
			// cons2
			multIn0aNext = MINUSONE; multIn0bNext = multOut0; 
			// m144
			multIn1aNext = reg713; multIn1bNext = TWO; 
			// m244
			multIn2aNext = reg714; multIn2bNext = TWO; 
			// d085
			divIn0aNext = reg442; divIn0bNext = reg447; 
			// a024
			reg444Next = addsubOut0;
			// cons1
			reg501Next = multOut0;
			// cons3
			reg648Next = multOut1;
			// cons4
			reg679Next = multOut2;
		end
		3:begin
			// a133
			addsubIn0aNext = reg444; addsubIn0bNext = addsubOut0; addsubMod0Next = add; 
			// s115
			addsubIn1aNext = reg113; addsubIn1bNext = divOut0; addsubMod1Next = sub; 
			if ( reg058 != 0 && reg025 == 0 ) begin
				addsubIn1aNext = ZERO; addsubIn1bNext = divOut0; addsubMod1Next = sub; 
			end
			// s276
			addsubIn2aNext = reg458; addsubIn2bNext = reg290; addsubMod2Next = sub; 
			// s393
			addsubIn3aNext = reg469; addsubIn3bNext = reg314; addsubMod3Next = sub; 
			// m004
			multIn0aNext = TAU; multIn0bNext = addsubOut2; 
			// m057
			multIn1aNext = reg715; multIn1bNext = TWO; 
			// cons6
			divIn0aNext = reg315; divIn0bNext = reg387; 
			// bool0
			eqgtgeltleneIn0aNext = addsubOut1; eqgtgeltleneIn0bNext = ONE; eqgtgeltleneMod0Next = lt; 
			// a035
			reg446Next = addsubOut1;
			// m283
			reg710Next = multOut0;
			// m382
			reg711Next = multOut1;
			// m482
			reg712Next = multOut2;
		end
		4:begin
			// s223
			addsubIn0aNext = reg162; addsubIn0bNext = divOut0; addsubMod0Next = sub; 
			if ( reg058 == 0 && reg025 != 0 ) begin
				addsubIn0aNext = ZERO; addsubIn0bNext = divOut0; addsubMod0Next = sub; 
			end
			// a158
			addsubIn1aNext = reg493; addsubIn1bNext = reg492; addsubMod1Next = add; 
			// a257
			addsubIn2aNext = reg386; addsubIn2bNext = reg490; addsubMod2Next = add; 
			// a374
			addsubIn3aNext = reg494; addsubIn3bNext = reg499; addsubMod3Next = add; 
			// m072
			multIn0aNext = addsubOut0; multIn0bNext = addsubOut0; 
			// m171
			multIn1aNext = addsubOut1; multIn1bNext = addsubOut1; 
			// m271
			multIn2aNext = addsubOut2; multIn2bNext = addsubOut2; 
			// cons7
			divIn0aNext = reg339; divIn0bNext = reg387; 
			// a062
			reg389Next = addsubOut0;
			// a161
			reg398Next = addsubOut1;
			// a261
			reg407Next = addsubOut2;
			// a322
			reg455Next = addsubOut3;
			// cons2
			reg531Next = multOut0;
			// m144
			reg716Next = multOut1;
			// m244
			reg717Next = multOut2;
		end
		5:begin
			// s058
			addsubIn0aNext = reg183; addsubIn0bNext = multOut0; addsubMod0Next = sub; 
			if ( reg064 == 0 && reg031 == 0 ) begin
				addsubIn0aNext = reg183; addsubIn0bNext = ZERO; addsubMod0Next = sub; 
			end
			// as335
			addsubIn1aNext = reg467; addsubIn1bNext = reg710; addsubMod1Next = sub; 
			if ( reg561 ) begin
				addsubIn1aNext = reg467; addsubIn1bNext = reg678; addsubMod1Next = sub; 
			end
			if ( reg563 ) begin
				addsubIn1aNext = reg467; addsubIn1bNext = reg678; addsubMod1Next = sub; 
			end
			// as432
			addsubIn2aNext = reg477; addsubIn2bNext = reg711; addsubMod2Next = sub; 
			if ( reg561 ) begin
				addsubIn2aNext = reg477; addsubIn2bNext = reg709; addsubMod2Next = sub; 
			end
			if ( reg563 ) begin
				addsubIn2aNext = reg477; addsubIn2bNext = reg709; addsubMod2Next = sub; 
			end
			// as049
			addsubIn3aNext = reg489; addsubIn3bNext = reg712; addsubMod3Next = sub; 
			if ( reg561 ) begin
				addsubIn3aNext = reg489; addsubIn3bNext = cons5; addsubMod3Next = sub; 
			end
			if ( reg563 ) begin
				addsubIn3aNext = reg489; addsubIn3bNext = cons5; addsubMod3Next = sub; 
			end
			// m371
			multIn0aNext = addsubOut0; multIn0bNext = addsubOut0; 
			// m471
			multIn1aNext = addsubOut1; multIn1bNext = addsubOut1; 
			// m083
			multIn2aNext = addsubOut2; multIn2bNext = addsubOut2; 
			// cons8
			divIn0aNext = reg388; divIn0bNext = reg387; 
			// ct1
			sqrtIn0aNext = reg445; 
			if ( eqgtgeltleneOut0 ) begin
				sqrtIn0aNext = ONE; 
			end
			// a361
			reg416Next = addsubOut0;
			// a461
			reg425Next = addsubOut1;
			// a073
			reg435Next = addsubOut2;
			// s171
			reg451Next = addsubOut3;
			// cons6
			reg564Next = divOut0;
			// m057
			reg718Next = multOut1;
		end
		6:begin
			// a024
			addsubIn0aNext = multOut1; addsubIn0bNext = multOut0; addsubMod0Next = add; 
			// s316
			addsubIn1aNext = reg716; addsubIn1bNext = reg197; addsubMod1Next = sub; 
			// s413
			addsubIn2aNext = reg717; addsubIn2bNext = reg232; addsubMod2Next = sub; 
			// s424
			addsubIn3aNext = reg718; addsubIn3bNext = reg267; addsubMod3Next = sub; 
			// m010
			multIn0aNext = carpan1; multIn0bNext = addsubOut0; 
			// m110
			multIn1aNext = carpan1; multIn1bNext = addsubOut1; 
			// m210
			multIn2aNext = carpan2; multIn2bNext = addsubOut2; 
			// s300
			reg415Next = addsubOut3;
			// m271
			reg443Next = multOut2;
			// c080
			reg560Next = eqgtgeltleneOut0;
			// cons7
			reg592Next = divOut0;
		end
		7:begin
			// a122
			addsubIn0aNext = multOut1; addsubIn0bNext = multOut0; addsubMod0Next = add; 
			// a035
			addsubIn1aNext = reg443; addsubIn1bNext = multOut2; addsubMod1Next = add; 
			// a196
			addsubIn2aNext = reg451; addsubIn2bNext = addsubOut3; addsubMod2Next = add; 
			// m310
			multIn0aNext = carpan1; multIn0bNext = reg415; 
			// m410
			multIn1aNext = carpan1; multIn1bNext = addsubOut0; 
			// m021
			multIn2aNext = carpan2; multIn2bNext = addsubOut1; 
			// d030
			divIn0aNext = reg397; divIn0bNext = sqrtOut0; 
			// ct1
			reg448Next = sqrtOut0;
			// s096
			reg452Next = addsubOut2;
			// c091
			reg562Next = eqgtgeltleneOut0;
			// cons8
			reg620Next = divOut0;
		end
		8:begin
			// a062
			addsubIn0aNext = reg004; addsubIn0bNext = multOut0; addsubMod0Next = add; 
			if ( reg013 == n ) begin
				addsubIn0aNext = ZERO; addsubIn0bNext = ZERO; addsubMod0Next = add; 
			end
			// a161
			addsubIn1aNext = reg007; addsubIn1bNext = multOut1; addsubMod1Next = add; 
			if ( reg013 == n ) begin
				addsubIn1aNext = ZERO; addsubIn1bNext = ZERO; addsubMod1Next = add; 
			end
			// a261
			addsubIn2aNext = reg010; addsubIn2bNext = multOut2; addsubMod2Next = add; 
			if ( reg013 == n ) begin
				addsubIn2aNext = ZERO; addsubIn2bNext = ZERO; addsubMod2Next = add; 
			end
			// a322
			addsubIn3aNext = reg452; addsubIn3bNext = addsubOut0; addsubMod3Next = add; 
			// m035
			multIn0aNext = TAU; multIn0bNext = reg455; 
			// m046
			multIn1aNext = TAU; multIn1bNext = addsubOut1; 
			// m202
			multIn2aNext = BETA; multIn2bNext = addsubOut3; 
			// d041
			divIn0aNext = reg406; divIn0bNext = reg448; 
			// s187
			reg468Next = addsubOut2;
			// s295
			reg478Next = addsubOut3;
		end
		9:begin
			// a361
			addsubIn0aNext = reg037; addsubIn0bNext = multOut0; addsubMod0Next = add; 
			if ( reg046 == m ) begin
				addsubIn0aNext = ZERO; addsubIn0bNext = ZERO; addsubMod0Next = add; 
			end
			// a461
			addsubIn1aNext = reg040; addsubIn1bNext = multOut1; addsubMod1Next = add; 
			if ( reg046 == m ) begin
				addsubIn1aNext = ZERO; addsubIn1bNext = ZERO; addsubMod1Next = add; 
			end
			// a073
			addsubIn2aNext = reg043; addsubIn2bNext = multOut2; addsubMod2Next = add; 
			if ( reg046 == m ) begin
				addsubIn2aNext = ZERO; addsubIn2bNext = ZERO; addsubMod2Next = add; 
			end
			// s171
			addsubIn3aNext = reg081; addsubIn3bNext = divOut0; addsubMod3Next = sub; 
			if ( reg059 != 0 && reg026 == 0 ) begin
				addsubIn3aNext = ZERO; addsubIn3bNext = divOut0; addsubMod3Next = sub; 
			end
			// m182
			multIn0aNext = addsubOut2; multIn0bNext = reg338; 
			// m103
			multIn1aNext = addsubOut3; multIn1bNext = reg363; 
			// d063
			divIn0aNext = reg424; divIn0bNext = reg448; 
			// ct0
			sqrtIn0aNext = reg446; 
			if ( eqgtgeltleneOut0 ) begin
				sqrtIn0aNext = ONE; 
			end
			// bool1
			eqgtgeltleneIn0aNext = addsubOut0; eqgtgeltleneIn0bNext = ONE; eqgtgeltleneMod0Next = lt; 
			// a133
			reg445Next = addsubOut0;
			// s115
			reg453Next = addsubOut1;
			reg390Next = reg389;
			reg391Next = reg390;
			reg392Next = reg391;
			reg393Next = reg392;
			reg394Next = reg393;
			reg395Next = reg394;
			reg396Next = reg395;
			reg397Next = reg396;
			reg399Next = reg398;
			reg400Next = reg399;
			reg401Next = reg400;
			reg402Next = reg401;
			reg403Next = reg402;
			reg404Next = reg403;
			reg405Next = reg404;
			reg406Next = reg405;
			reg408Next = reg407;
			reg409Next = reg408;
			reg410Next = reg409;
			reg411Next = reg410;
			reg412Next = reg411;
			reg413Next = reg412;
			reg414Next = reg413;
			reg417Next = reg416;
			reg418Next = reg417;
			reg419Next = reg418;
			reg420Next = reg419;
			reg421Next = reg420;
			reg422Next = reg421;
			reg423Next = reg422;
			reg424Next = reg423;
			reg426Next = reg425;
			reg427Next = reg426;
			reg428Next = reg427;
			reg429Next = reg428;
			reg430Next = reg429;
			reg431Next = reg430;
			reg432Next = reg431;
			reg433Next = reg432;
			reg434Next = reg433;
			reg436Next = reg435;
			reg437Next = reg436;
			reg438Next = reg437;
			reg439Next = reg438;
			reg440Next = reg439;
			reg441Next = reg440;
			reg442Next = reg441;
			reg449Next = reg448;
			reg459Next = reg458;
			reg460Next = reg459;
			reg461Next = reg460;
			reg462Next = reg461;
			reg463Next = reg462;
			reg464Next = reg463;
			reg465Next = reg464;
			reg466Next = reg465;
			reg467Next = reg466;
			reg469Next = reg468;
			reg470Next = reg469;
			reg471Next = reg470;
			reg472Next = reg471;
			reg473Next = reg472;
			reg474Next = reg473;
			reg475Next = reg474;
			reg476Next = reg475;
			reg477Next = reg476;
			reg479Next = reg478;
			reg480Next = reg479;
			reg481Next = reg480;
			reg482Next = reg481;
			reg483Next = reg482;
			reg484Next = reg483;
			reg485Next = reg484;
			reg486Next = reg485;
			reg487Next = reg486;
			reg488Next = reg487;
			reg489Next = reg488;
			reg492Next = reg491;
			reg496Next = reg495;
			reg497Next = reg496;
			reg498Next = reg497;
			reg499Next = reg498;
			reg502Next = reg501;
			reg503Next = reg502;
			reg504Next = reg503;
			reg505Next = reg504;
			reg506Next = reg505;
			reg507Next = reg506;
			reg508Next = reg507;
			reg509Next = reg508;
			reg510Next = reg509;
			reg511Next = reg510;
			reg512Next = reg511;
			reg513Next = reg512;
			reg514Next = reg513;
			reg515Next = reg514;
			reg516Next = reg515;
			reg517Next = reg516;
			reg518Next = reg517;
			reg519Next = reg518;
			reg520Next = reg519;
			reg521Next = reg520;
			reg522Next = reg521;
			reg523Next = reg522;
			reg524Next = reg523;
			reg525Next = reg524;
			reg526Next = reg525;
			reg527Next = reg526;
			reg528Next = reg527;
			reg529Next = reg528;
			reg530Next = reg529;
			reg532Next = reg531;
			reg533Next = reg532;
			reg534Next = reg533;
			reg535Next = reg534;
			reg536Next = reg535;
			reg537Next = reg536;
			reg538Next = reg537;
			reg539Next = reg538;
			reg540Next = reg539;
			reg541Next = reg540;
			reg542Next = reg541;
			reg543Next = reg542;
			reg544Next = reg543;
			reg545Next = reg544;
			reg546Next = reg545;
			reg547Next = reg546;
			reg548Next = reg547;
			reg549Next = reg548;
			reg550Next = reg549;
			reg551Next = reg550;
			reg552Next = reg551;
			reg553Next = reg552;
			reg554Next = reg553;
			reg555Next = reg554;
			reg556Next = reg555;
			reg557Next = reg556;
			reg558Next = reg557;
			reg559Next = reg558;
			reg561Next = reg560;
			reg563Next = reg562;
			reg565Next = reg564;
			reg566Next = reg565;
			reg567Next = reg566;
			reg568Next = reg567;
			reg569Next = reg568;
			reg570Next = reg569;
			reg571Next = reg570;
			reg572Next = reg571;
			reg573Next = reg572;
			reg574Next = reg573;
			reg575Next = reg574;
			reg576Next = reg575;
			reg577Next = reg576;
			reg578Next = reg577;
			reg579Next = reg578;
			reg580Next = reg579;
			reg581Next = reg580;
			reg582Next = reg581;
			reg583Next = reg582;
			reg584Next = reg583;
			reg585Next = reg584;
			reg586Next = reg585;
			reg587Next = reg586;
			reg588Next = reg587;
			reg589Next = reg588;
			reg590Next = reg589;
			reg591Next = reg590;
			reg593Next = reg592;
			reg594Next = reg593;
			reg595Next = reg594;
			reg596Next = reg595;
			reg597Next = reg596;
			reg598Next = reg597;
			reg599Next = reg598;
			reg600Next = reg599;
			reg601Next = reg600;
			reg602Next = reg601;
			reg603Next = reg602;
			reg604Next = reg603;
			reg605Next = reg604;
			reg606Next = reg605;
			reg607Next = reg606;
			reg608Next = reg607;
			reg609Next = reg608;
			reg610Next = reg609;
			reg611Next = reg610;
			reg612Next = reg611;
			reg613Next = reg612;
			reg614Next = reg613;
			reg615Next = reg614;
			reg616Next = reg615;
			reg617Next = reg616;
			reg618Next = reg617;
			reg619Next = reg618;
			reg621Next = reg620;
			reg622Next = reg621;
			reg623Next = reg622;
			reg624Next = reg623;
			reg625Next = reg624;
			reg626Next = reg625;
			reg627Next = reg626;
			reg628Next = reg627;
			reg629Next = reg628;
			reg630Next = reg629;
			reg631Next = reg630;
			reg632Next = reg631;
			reg633Next = reg632;
			reg634Next = reg633;
			reg635Next = reg634;
			reg636Next = reg635;
			reg637Next = reg636;
			reg638Next = reg637;
			reg639Next = reg638;
			reg640Next = reg639;
			reg641Next = reg640;
			reg642Next = reg641;
			reg643Next = reg642;
			reg644Next = reg643;
			reg645Next = reg644;
			reg646Next = reg645;
			reg647Next = reg646;
			reg649Next = reg648;
			reg650Next = reg649;
			reg651Next = reg650;
			reg652Next = reg651;
			reg653Next = reg652;
			reg654Next = reg653;
			reg655Next = reg654;
			reg656Next = reg655;
			reg657Next = reg656;
			reg658Next = reg657;
			reg659Next = reg658;
			reg660Next = reg659;
			reg661Next = reg660;
			reg662Next = reg661;
			reg663Next = reg662;
			reg664Next = reg663;
			reg665Next = reg664;
			reg666Next = reg665;
			reg667Next = reg666;
			reg668Next = reg667;
			reg669Next = reg668;
			reg670Next = reg669;
			reg671Next = reg670;
			reg672Next = reg671;
			reg673Next = reg672;
			reg674Next = reg673;
			reg675Next = reg674;
			reg676Next = reg675;
			reg677Next = reg676;
			reg678Next = reg677;
			reg680Next = reg679;
			reg681Next = reg680;
			reg682Next = reg681;
			reg683Next = reg682;
			reg684Next = reg683;
			reg685Next = reg684;
			reg686Next = reg685;
			reg687Next = reg686;
			reg688Next = reg687;
			reg689Next = reg688;
			reg690Next = reg689;
			reg691Next = reg690;
			reg692Next = reg691;
			reg693Next = reg692;
			reg694Next = reg693;
			reg695Next = reg694;
			reg696Next = reg695;
			reg697Next = reg696;
			reg698Next = reg697;
			reg699Next = reg698;
			reg700Next = reg699;
			reg701Next = reg700;
			reg702Next = reg701;
			reg703Next = reg702;
			reg704Next = reg703;
			reg705Next = reg704;
			reg706Next = reg705;
			reg707Next = reg706;
			reg708Next = reg707;
			reg709Next = reg708;
			reg003Next = reg002;
			reg004Next = reg003;
			reg006Next = reg005;
			reg007Next = reg006;
			reg009Next = reg008;
			reg010Next = reg009;
			reg012Next = reg011;
			reg013Next = reg012;
			reg014Next = reg013;
			reg015Next = reg014;
			reg016Next = reg015;
			reg017Next = reg016;
			reg018Next = reg017;
			reg019Next = reg018;
			reg020Next = reg019;
			reg021Next = reg020;
			reg022Next = reg021;
			reg023Next = reg022;
			reg024Next = reg023;
			reg025Next = reg024;
			reg026Next = reg025;
			reg027Next = reg026;
			reg028Next = reg027;
			reg029Next = reg028;
			reg030Next = reg029;
			reg031Next = reg030;
			reg032Next = reg031;
			reg036Next = reg035;
			reg037Next = reg036;
			reg039Next = reg038;
			reg040Next = reg039;
			reg042Next = reg041;
			reg043Next = reg042;
			reg045Next = reg044;
			reg046Next = reg045;
			reg047Next = reg046;
			reg048Next = reg047;
			reg049Next = reg048;
			reg050Next = reg049;
			reg051Next = reg050;
			reg052Next = reg051;
			reg053Next = reg052;
			reg054Next = reg053;
			reg055Next = reg054;
			reg056Next = reg055;
			reg057Next = reg056;
			reg058Next = reg057;
			reg059Next = reg058;
			reg060Next = reg059;
			reg061Next = reg060;
			reg062Next = reg061;
			reg063Next = reg062;
			reg064Next = reg063;
			reg065Next = reg064;
			reg067Next = reg066;
			reg068Next = reg067;
			reg069Next = reg068;
			reg070Next = reg069;
			reg071Next = reg070;
			reg072Next = reg071;
			reg073Next = reg072;
			reg074Next = reg073;
			reg075Next = reg074;
			reg076Next = reg075;
			reg077Next = reg076;
			reg078Next = reg077;
			reg079Next = reg078;
			reg080Next = reg079;
			reg081Next = reg080;
			reg083Next = reg082;
			reg084Next = reg083;
			reg085Next = reg084;
			reg086Next = reg085;
			reg087Next = reg086;
			reg088Next = reg087;
			reg089Next = reg088;
			reg090Next = reg089;
			reg091Next = reg090;
			reg092Next = reg091;
			reg093Next = reg092;
			reg094Next = reg093;
			reg095Next = reg094;
			reg096Next = reg095;
			reg097Next = reg096;
			reg098Next = reg097;
			reg100Next = reg099;
			reg101Next = reg100;
			reg102Next = reg101;
			reg103Next = reg102;
			reg104Next = reg103;
			reg105Next = reg104;
			reg106Next = reg105;
			reg107Next = reg106;
			reg108Next = reg107;
			reg109Next = reg108;
			reg110Next = reg109;
			reg111Next = reg110;
			reg112Next = reg111;
			reg113Next = reg112;
			reg115Next = reg114;
			reg116Next = reg115;
			reg117Next = reg116;
			reg118Next = reg117;
			reg119Next = reg118;
			reg120Next = reg119;
			reg121Next = reg120;
			reg122Next = reg121;
			reg123Next = reg122;
			reg124Next = reg123;
			reg125Next = reg124;
			reg126Next = reg125;
			reg127Next = reg126;
			reg128Next = reg127;
			reg129Next = reg128;
			reg130Next = reg129;
			reg132Next = reg131;
			reg133Next = reg132;
			reg134Next = reg133;
			reg135Next = reg134;
			reg136Next = reg135;
			reg137Next = reg136;
			reg138Next = reg137;
			reg139Next = reg138;
			reg140Next = reg139;
			reg141Next = reg140;
			reg142Next = reg141;
			reg143Next = reg142;
			reg144Next = reg143;
			reg145Next = reg144;
			reg146Next = reg145;
			reg147Next = reg146;
			reg149Next = reg148;
			reg150Next = reg149;
			reg151Next = reg150;
			reg152Next = reg151;
			reg153Next = reg152;
			reg154Next = reg153;
			reg155Next = reg154;
			reg156Next = reg155;
			reg157Next = reg156;
			reg158Next = reg157;
			reg159Next = reg158;
			reg160Next = reg159;
			reg161Next = reg160;
			reg162Next = reg161;
			reg164Next = reg163;
			reg165Next = reg164;
			reg166Next = reg165;
			reg167Next = reg166;
			reg168Next = reg167;
			reg169Next = reg168;
			reg170Next = reg169;
			reg171Next = reg170;
			reg172Next = reg171;
			reg173Next = reg172;
			reg174Next = reg173;
			reg175Next = reg174;
			reg176Next = reg175;
			reg177Next = reg176;
			reg178Next = reg177;
			reg179Next = reg178;
			reg180Next = reg179;
			reg181Next = reg180;
			reg182Next = reg181;
			reg183Next = reg182;
			reg184Next = reg183;
			reg185Next = reg184;
			reg186Next = reg185;
			reg187Next = reg186;
			reg188Next = reg187;
			reg189Next = reg188;
			reg190Next = reg189;
			reg191Next = reg190;
			reg192Next = reg191;
			reg193Next = reg192;
			reg194Next = reg193;
			reg195Next = reg194;
			reg196Next = reg195;
			reg197Next = reg196;
			reg199Next = reg198;
			reg200Next = reg199;
			reg201Next = reg200;
			reg202Next = reg201;
			reg203Next = reg202;
			reg204Next = reg203;
			reg205Next = reg204;
			reg206Next = reg205;
			reg207Next = reg206;
			reg208Next = reg207;
			reg209Next = reg208;
			reg210Next = reg209;
			reg211Next = reg210;
			reg212Next = reg211;
			reg213Next = reg212;
			reg214Next = reg213;
			reg215Next = reg214;
			reg216Next = reg215;
			reg217Next = reg216;
			reg218Next = reg217;
			reg219Next = reg218;
			reg220Next = reg219;
			reg221Next = reg220;
			reg222Next = reg221;
			reg223Next = reg222;
			reg224Next = reg223;
			reg225Next = reg224;
			reg226Next = reg225;
			reg227Next = reg226;
			reg228Next = reg227;
			reg229Next = reg228;
			reg230Next = reg229;
			reg231Next = reg230;
			reg232Next = reg231;
			reg234Next = reg233;
			reg235Next = reg234;
			reg236Next = reg235;
			reg237Next = reg236;
			reg238Next = reg237;
			reg239Next = reg238;
			reg240Next = reg239;
			reg241Next = reg240;
			reg242Next = reg241;
			reg243Next = reg242;
			reg244Next = reg243;
			reg245Next = reg244;
			reg246Next = reg245;
			reg247Next = reg246;
			reg248Next = reg247;
			reg249Next = reg248;
			reg250Next = reg249;
			reg251Next = reg250;
			reg252Next = reg251;
			reg253Next = reg252;
			reg254Next = reg253;
			reg255Next = reg254;
			reg256Next = reg255;
			reg257Next = reg256;
			reg258Next = reg257;
			reg259Next = reg258;
			reg260Next = reg259;
			reg261Next = reg260;
			reg262Next = reg261;
			reg263Next = reg262;
			reg264Next = reg263;
			reg265Next = reg264;
			reg266Next = reg265;
			reg267Next = reg266;
			reg269Next = reg268;
			reg270Next = reg269;
			reg271Next = reg270;
			reg272Next = reg271;
			reg273Next = reg272;
			reg274Next = reg273;
			reg275Next = reg274;
			reg276Next = reg275;
			reg277Next = reg276;
			reg278Next = reg277;
			reg279Next = reg278;
			reg280Next = reg279;
			reg281Next = reg280;
			reg282Next = reg281;
			reg283Next = reg282;
			reg284Next = reg283;
			reg285Next = reg284;
			reg286Next = reg285;
			reg287Next = reg286;
			reg288Next = reg287;
			reg289Next = reg288;
			reg290Next = reg289;
			reg292Next = reg291;
			reg293Next = reg292;
			reg294Next = reg293;
			reg295Next = reg294;
			reg296Next = reg295;
			reg297Next = reg296;
			reg298Next = reg297;
			reg299Next = reg298;
			reg300Next = reg299;
			reg301Next = reg300;
			reg302Next = reg301;
			reg303Next = reg302;
			reg304Next = reg303;
			reg305Next = reg304;
			reg306Next = reg305;
			reg307Next = reg306;
			reg308Next = reg307;
			reg309Next = reg308;
			reg310Next = reg309;
			reg311Next = reg310;
			reg312Next = reg311;
			reg313Next = reg312;
			reg314Next = reg313;
			reg316Next = reg315;
			reg317Next = reg316;
			reg318Next = reg317;
			reg319Next = reg318;
			reg320Next = reg319;
			reg321Next = reg320;
			reg322Next = reg321;
			reg323Next = reg322;
			reg324Next = reg323;
			reg325Next = reg324;
			reg326Next = reg325;
			reg327Next = reg326;
			reg328Next = reg327;
			reg329Next = reg328;
			reg330Next = reg329;
			reg331Next = reg330;
			reg332Next = reg331;
			reg333Next = reg332;
			reg334Next = reg333;
			reg335Next = reg334;
			reg336Next = reg335;
			reg337Next = reg336;
			reg338Next = reg337;
			reg340Next = reg339;
			reg341Next = reg340;
			reg342Next = reg341;
			reg343Next = reg342;
			reg344Next = reg343;
			reg345Next = reg344;
			reg346Next = reg345;
			reg347Next = reg346;
			reg348Next = reg347;
			reg349Next = reg348;
			reg350Next = reg349;
			reg351Next = reg350;
			reg352Next = reg351;
			reg353Next = reg352;
			reg354Next = reg353;
			reg355Next = reg354;
			reg356Next = reg355;
			reg357Next = reg356;
			reg358Next = reg357;
			reg359Next = reg358;
			reg360Next = reg359;
			reg361Next = reg360;
			reg362Next = reg361;
			reg363Next = reg362;
			reg365Next = reg364;
			reg366Next = reg365;
			reg367Next = reg366;
			reg368Next = reg367;
			reg369Next = reg368;
			reg370Next = reg369;
			reg371Next = reg370;
			reg372Next = reg371;
			reg373Next = reg372;
			reg374Next = reg373;
			reg375Next = reg374;
			reg376Next = reg375;
			reg377Next = reg376;
			reg378Next = reg377;
			reg379Next = reg378;
			reg380Next = reg379;
			reg381Next = reg380;
			reg382Next = reg381;
			reg383Next = reg382;
			reg384Next = reg383;
			reg385Next = reg384;
			reg386Next = reg385;
		end
		default: begin
		end
		endcase
	end
endmodule
